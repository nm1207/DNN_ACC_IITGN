// This is the unpowered netlist.
module mac (clk,
    reset,
    data_in,
    data_out);
 input clk;
 input reset;
 input [255:0] data_in;
 output [27:0] data_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net113));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_4 _06438_ (.A(net257),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_4 _06439_ (.A(_02174_),
    .X(_02185_));
 sky130_fd_sc_hd__clkbuf_4 _06440_ (.A(net24),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_4 _06441_ (.A(net15),
    .X(_02207_));
 sky130_fd_sc_hd__clkbuf_4 _06442_ (.A(net130),
    .X(_02218_));
 sky130_fd_sc_hd__buf_4 _06443_ (.A(net121),
    .X(_02229_));
 sky130_fd_sc_hd__buf_4 _06444_ (.A(net94),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_4 _06445_ (.A(net85),
    .X(_02251_));
 sky130_fd_sc_hd__a22o_1 _06446_ (.A1(_02218_),
    .A2(_02229_),
    .B1(_02240_),
    .B2(_02251_),
    .X(_02262_));
 sky130_fd_sc_hd__and4_2 _06447_ (.A(_02218_),
    .B(_02229_),
    .C(_02240_),
    .D(_02251_),
    .X(_02273_));
 sky130_fd_sc_hd__inv_2 _06448_ (.A(_02273_),
    .Y(_02284_));
 sky130_fd_sc_hd__nand4_2 _06449_ (.A(_02196_),
    .B(_02207_),
    .C(_02262_),
    .D(_02284_),
    .Y(_02295_));
 sky130_fd_sc_hd__a22o_1 _06450_ (.A1(_02196_),
    .A2(_02207_),
    .B1(_02262_),
    .B2(_02284_),
    .X(_02306_));
 sky130_fd_sc_hd__buf_2 _06451_ (.A(net165),
    .X(_02317_));
 sky130_fd_sc_hd__buf_2 _06452_ (.A(net157),
    .X(_02328_));
 sky130_fd_sc_hd__and2_1 _06453_ (.A(_02317_),
    .B(_02328_),
    .X(_02339_));
 sky130_fd_sc_hd__and3_2 _06454_ (.A(_02295_),
    .B(_02306_),
    .C(_02339_),
    .X(_02350_));
 sky130_fd_sc_hd__a21oi_1 _06455_ (.A1(_02295_),
    .A2(_02306_),
    .B1(_02339_),
    .Y(_02361_));
 sky130_fd_sc_hd__or2_1 _06456_ (.A(_02350_),
    .B(_02361_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_4 _06457_ (.A(net148),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_4 _06458_ (.A(net139),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_2 _06459_ (.A(_02383_),
    .B(_02394_),
    .Y(_02405_));
 sky130_fd_sc_hd__or2_1 _06460_ (.A(_02372_),
    .B(_02405_),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_1 _06461_ (.A(_02372_),
    .B(_02405_),
    .Y(_02426_));
 sky130_fd_sc_hd__and2_1 _06462_ (.A(_02415_),
    .B(_02426_),
    .X(_02437_));
 sky130_fd_sc_hd__clkbuf_4 _06463_ (.A(net208),
    .X(_02448_));
 sky130_fd_sc_hd__clkbuf_4 _06464_ (.A(net199),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_4 _06465_ (.A(net6),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_4 _06466_ (.A(net252),
    .X(_02481_));
 sky130_fd_sc_hd__buf_4 _06467_ (.A(net243),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_4 _06468_ (.A(net235),
    .X(_02503_));
 sky130_fd_sc_hd__a22o_1 _06469_ (.A1(_02470_),
    .A2(_02481_),
    .B1(_02492_),
    .B2(_02503_),
    .X(_02514_));
 sky130_fd_sc_hd__nand4_4 _06470_ (.A(_02470_),
    .B(_02481_),
    .C(_02492_),
    .D(_02503_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand4_4 _06471_ (.A(_02448_),
    .B(_02459_),
    .C(_02514_),
    .D(_02525_),
    .Y(_02536_));
 sky130_fd_sc_hd__a22o_2 _06472_ (.A1(_02448_),
    .A2(_02459_),
    .B1(_02514_),
    .B2(_02525_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _06473_ (.A(_02536_),
    .B(_02547_),
    .Y(_02558_));
 sky130_fd_sc_hd__clkbuf_4 _06474_ (.A(net59),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_4 _06475_ (.A(net50),
    .X(_02580_));
 sky130_fd_sc_hd__nand2_2 _06476_ (.A(_02569_),
    .B(_02580_),
    .Y(_02591_));
 sky130_fd_sc_hd__or2_1 _06477_ (.A(_02558_),
    .B(_02591_),
    .X(_02602_));
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(_02558_),
    .B(_02591_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(_02602_),
    .B(_02613_),
    .Y(_02624_));
 sky130_fd_sc_hd__buf_2 _06480_ (.A(net113),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_4 _06481_ (.A(net103),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_4 _06482_ (.A(net76),
    .X(_02657_));
 sky130_fd_sc_hd__buf_2 _06483_ (.A(net68),
    .X(_02668_));
 sky130_fd_sc_hd__a22o_1 _06484_ (.A1(_02635_),
    .A2(_02646_),
    .B1(_02657_),
    .B2(_02668_),
    .X(_02679_));
 sky130_fd_sc_hd__inv_2 _06485_ (.A(_02679_),
    .Y(_02690_));
 sky130_fd_sc_hd__and4_1 _06486_ (.A(_02635_),
    .B(_02646_),
    .C(_02657_),
    .D(_02668_),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_4 _06487_ (.A(net191),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_4 _06488_ (.A(net182),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_4 _06489_ (.A(net167),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_4 _06490_ (.A(net78),
    .X(_02745_));
 sky130_fd_sc_hd__a22oi_1 _06491_ (.A1(_02712_),
    .A2(_02723_),
    .B1(_02734_),
    .B2(_02745_),
    .Y(_02756_));
 sky130_fd_sc_hd__and4_1 _06492_ (.A(_02712_),
    .B(_02723_),
    .C(_02734_),
    .D(_02745_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _06493_ (.A(_02756_),
    .B(_02767_),
    .Y(_02778_));
 sky130_fd_sc_hd__buf_6 _06494_ (.A(net245),
    .X(_02789_));
 sky130_fd_sc_hd__clkbuf_4 _06495_ (.A(net1),
    .X(_02800_));
 sky130_fd_sc_hd__buf_4 _06496_ (.A(net41),
    .X(_02811_));
 sky130_fd_sc_hd__buf_4 _06497_ (.A(net32),
    .X(_02822_));
 sky130_fd_sc_hd__a22oi_4 _06498_ (.A1(_02789_),
    .A2(_02800_),
    .B1(_02811_),
    .B2(_02822_),
    .Y(_02833_));
 sky130_fd_sc_hd__and4_4 _06499_ (.A(_02789_),
    .B(_02800_),
    .C(_02811_),
    .D(_02822_),
    .X(_02844_));
 sky130_fd_sc_hd__buf_2 _06500_ (.A(net226),
    .X(_02855_));
 sky130_fd_sc_hd__buf_2 _06501_ (.A(net217),
    .X(_02866_));
 sky130_fd_sc_hd__or4bb_2 _06502_ (.A(_02833_),
    .B(_02844_),
    .C_N(_02855_),
    .D_N(_02866_),
    .X(_02877_));
 sky130_fd_sc_hd__a2bb2o_1 _06503_ (.A1_N(_02833_),
    .A2_N(_02844_),
    .B1(_02855_),
    .B2(_02866_),
    .X(_02888_));
 sky130_fd_sc_hd__and3_2 _06504_ (.A(_02778_),
    .B(_02877_),
    .C(_02888_),
    .X(_02899_));
 sky130_fd_sc_hd__and2_1 _06505_ (.A(_02877_),
    .B(_02888_),
    .X(_02910_));
 sky130_fd_sc_hd__nor2_1 _06506_ (.A(_02778_),
    .B(_02910_),
    .Y(_02921_));
 sky130_fd_sc_hd__or2_1 _06507_ (.A(_02899_),
    .B(_02921_),
    .X(_02932_));
 sky130_fd_sc_hd__nor3_1 _06508_ (.A(_02690_),
    .B(_02701_),
    .C(_02932_),
    .Y(_02943_));
 sky130_fd_sc_hd__o21a_1 _06509_ (.A1(_02690_),
    .A2(_02701_),
    .B1(_02932_),
    .X(_02954_));
 sky130_fd_sc_hd__or2_1 _06510_ (.A(_02943_),
    .B(_02954_),
    .X(_02965_));
 sky130_fd_sc_hd__nor2_1 _06511_ (.A(_02624_),
    .B(_02965_),
    .Y(_02976_));
 sky130_fd_sc_hd__inv_2 _06512_ (.A(_02976_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand2_1 _06513_ (.A(_02624_),
    .B(_02965_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand3_2 _06514_ (.A(_02437_),
    .B(_02987_),
    .C(_02998_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21o_1 _06515_ (.A1(_02987_),
    .A2(_02998_),
    .B1(_02437_),
    .X(_03020_));
 sky130_fd_sc_hd__a21o_1 _06516_ (.A1(_03009_),
    .A2(_03020_),
    .B1(net258),
    .X(_03031_));
 sky130_fd_sc_hd__nand3_1 _06517_ (.A(net258),
    .B(_03009_),
    .C(_03020_),
    .Y(_03042_));
 sky130_fd_sc_hd__and3_1 _06518_ (.A(_02185_),
    .B(_03031_),
    .C(_03042_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _06519_ (.A(_03053_),
    .X(_00000_));
 sky130_fd_sc_hd__and3_1 _06520_ (.A(_02437_),
    .B(_02987_),
    .C(_02998_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_4 _06521_ (.A(net33),
    .X(_03084_));
 sky130_fd_sc_hd__buf_2 _06522_ (.A(net112),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_4 _06523_ (.A(net256),
    .X(_03106_));
 sky130_fd_sc_hd__a22o_1 _06524_ (.A1(_03095_),
    .A2(_02789_),
    .B1(_03106_),
    .B2(_02800_),
    .X(_03117_));
 sky130_fd_sc_hd__and3_4 _06525_ (.A(net112),
    .B(net245),
    .C(net256),
    .X(_03128_));
 sky130_fd_sc_hd__nand2_4 _06526_ (.A(_02800_),
    .B(_03128_),
    .Y(_03139_));
 sky130_fd_sc_hd__and4_2 _06527_ (.A(net41),
    .B(_03084_),
    .C(_03117_),
    .D(_03139_),
    .X(_03150_));
 sky130_fd_sc_hd__a22oi_2 _06528_ (.A1(net41),
    .A2(_03084_),
    .B1(_03117_),
    .B2(_03139_),
    .Y(_03161_));
 sky130_fd_sc_hd__nor2_2 _06529_ (.A(_03150_),
    .B(_03161_),
    .Y(_03172_));
 sky130_fd_sc_hd__xor2_4 _06530_ (.A(_02844_),
    .B(_03172_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_4 _06531_ (.A(net42),
    .X(_03194_));
 sky130_fd_sc_hd__nand2_2 _06532_ (.A(_02822_),
    .B(_03194_),
    .Y(_03205_));
 sky130_fd_sc_hd__xnor2_4 _06533_ (.A(_03183_),
    .B(_03205_),
    .Y(_03216_));
 sky130_fd_sc_hd__buf_2 _06534_ (.A(net218),
    .X(_03227_));
 sky130_fd_sc_hd__and3_1 _06535_ (.A(_03227_),
    .B(net226),
    .C(net227),
    .X(_03238_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(_02866_),
    .B(_03238_),
    .Y(_03249_));
 sky130_fd_sc_hd__buf_2 _06537_ (.A(net227),
    .X(_03260_));
 sky130_fd_sc_hd__a22o_1 _06538_ (.A1(_03227_),
    .A2(_02855_),
    .B1(_03260_),
    .B2(_02866_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2_1 _06539_ (.A(_03249_),
    .B(_03271_),
    .Y(_03282_));
 sky130_fd_sc_hd__xor2_2 _06540_ (.A(_03216_),
    .B(_03282_),
    .X(_03293_));
 sky130_fd_sc_hd__or2_1 _06541_ (.A(_02877_),
    .B(_03293_),
    .X(_03304_));
 sky130_fd_sc_hd__nand2_1 _06542_ (.A(_02877_),
    .B(_03293_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(_03304_),
    .B(_03315_),
    .Y(_03326_));
 sky130_fd_sc_hd__clkbuf_4 _06544_ (.A(net183),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_4 _06545_ (.A(net192),
    .X(_03348_));
 sky130_fd_sc_hd__a22o_1 _06546_ (.A1(_03337_),
    .A2(_02712_),
    .B1(_03348_),
    .B2(_02723_),
    .X(_03359_));
 sky130_fd_sc_hd__nand4_1 _06547_ (.A(_03337_),
    .B(_02712_),
    .C(_03348_),
    .D(_02723_),
    .Y(_03370_));
 sky130_fd_sc_hd__clkbuf_4 _06548_ (.A(net89),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_4 _06549_ (.A(net174),
    .X(_03392_));
 sky130_fd_sc_hd__a22o_1 _06550_ (.A1(_03381_),
    .A2(_02734_),
    .B1(_03392_),
    .B2(_02745_),
    .X(_03403_));
 sky130_fd_sc_hd__and4_1 _06551_ (.A(_03381_),
    .B(net167),
    .C(_03392_),
    .D(_02745_),
    .X(_03414_));
 sky130_fd_sc_hd__inv_2 _06552_ (.A(_03414_),
    .Y(_03425_));
 sky130_fd_sc_hd__and4_1 _06553_ (.A(_03359_),
    .B(_03370_),
    .C(_03403_),
    .D(_03425_),
    .X(_03436_));
 sky130_fd_sc_hd__a22oi_1 _06554_ (.A1(_03359_),
    .A2(_03370_),
    .B1(_03403_),
    .B2(_03425_),
    .Y(_03447_));
 sky130_fd_sc_hd__nor2_1 _06555_ (.A(_03436_),
    .B(_03447_),
    .Y(_03458_));
 sky130_fd_sc_hd__and2_1 _06556_ (.A(_02767_),
    .B(_03458_),
    .X(_03469_));
 sky130_fd_sc_hd__nor2_1 _06557_ (.A(_02767_),
    .B(_03458_),
    .Y(_03480_));
 sky130_fd_sc_hd__or2_1 _06558_ (.A(_03469_),
    .B(_03480_),
    .X(_03491_));
 sky130_fd_sc_hd__xor2_2 _06559_ (.A(_03326_),
    .B(_03491_),
    .X(_03502_));
 sky130_fd_sc_hd__xnor2_1 _06560_ (.A(_02899_),
    .B(_03502_),
    .Y(_03513_));
 sky130_fd_sc_hd__clkbuf_4 _06561_ (.A(net104),
    .X(_03524_));
 sky130_fd_sc_hd__and3_1 _06562_ (.A(_03524_),
    .B(net113),
    .C(net114),
    .X(_03535_));
 sky130_fd_sc_hd__buf_2 _06563_ (.A(net114),
    .X(_03546_));
 sky130_fd_sc_hd__a22o_1 _06564_ (.A1(_03524_),
    .A2(_02635_),
    .B1(_03546_),
    .B2(_02646_),
    .X(_03557_));
 sky130_fd_sc_hd__a21bo_1 _06565_ (.A1(_02646_),
    .A2(_03535_),
    .B1_N(_03557_),
    .X(_03568_));
 sky130_fd_sc_hd__buf_2 _06566_ (.A(net69),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_4 _06567_ (.A(net77),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_1 _06568_ (.A1(_03579_),
    .A2(_02657_),
    .B1(_03590_),
    .B2(_02668_),
    .X(_03601_));
 sky130_fd_sc_hd__and3_1 _06569_ (.A(_03579_),
    .B(_02657_),
    .C(_03590_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(_02668_),
    .B(_03612_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(_03601_),
    .B(_03623_),
    .Y(_03634_));
 sky130_fd_sc_hd__xor2_1 _06572_ (.A(_03568_),
    .B(_03634_),
    .X(_03645_));
 sky130_fd_sc_hd__and2_1 _06573_ (.A(_02701_),
    .B(_03645_),
    .X(_03656_));
 sky130_fd_sc_hd__nor2_1 _06574_ (.A(_02701_),
    .B(_03645_),
    .Y(_03667_));
 sky130_fd_sc_hd__or2_1 _06575_ (.A(_03656_),
    .B(_03667_),
    .X(_03678_));
 sky130_fd_sc_hd__or2_1 _06576_ (.A(_03513_),
    .B(_03678_),
    .X(_03689_));
 sky130_fd_sc_hd__nand2_1 _06577_ (.A(_03513_),
    .B(_03678_),
    .Y(_03699_));
 sky130_fd_sc_hd__nand3_1 _06578_ (.A(_02943_),
    .B(_03689_),
    .C(_03699_),
    .Y(_03710_));
 sky130_fd_sc_hd__a21o_1 _06579_ (.A1(_03689_),
    .A2(_03699_),
    .B1(_02943_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_4 _06580_ (.A(net51),
    .X(_03732_));
 sky130_fd_sc_hd__buf_2 _06581_ (.A(net60),
    .X(_03743_));
 sky130_fd_sc_hd__a22oi_1 _06582_ (.A1(_03732_),
    .A2(_02569_),
    .B1(_03743_),
    .B2(_02580_),
    .Y(_03754_));
 sky130_fd_sc_hd__and4_1 _06583_ (.A(_03732_),
    .B(_02569_),
    .C(_03743_),
    .D(_02580_),
    .X(_03765_));
 sky130_fd_sc_hd__nor2_1 _06584_ (.A(_03754_),
    .B(_03765_),
    .Y(_03776_));
 sky130_fd_sc_hd__and3_1 _06585_ (.A(net253),
    .B(net6),
    .C(net7),
    .X(_03787_));
 sky130_fd_sc_hd__buf_2 _06586_ (.A(net7),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_1 _06587_ (.A(_03798_),
    .B(_02481_),
    .Y(_03809_));
 sky130_fd_sc_hd__clkbuf_4 _06588_ (.A(net253),
    .X(_03820_));
 sky130_fd_sc_hd__nand2_1 _06589_ (.A(_03820_),
    .B(_02470_),
    .Y(_03831_));
 sky130_fd_sc_hd__a22o_2 _06590_ (.A1(_02481_),
    .A2(_03787_),
    .B1(_03809_),
    .B2(_03831_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_4 _06591_ (.A(net236),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_4 _06592_ (.A(net244),
    .X(_03864_));
 sky130_fd_sc_hd__a22o_1 _06593_ (.A1(_03853_),
    .A2(_02492_),
    .B1(_03864_),
    .B2(_02503_),
    .X(_03875_));
 sky130_fd_sc_hd__and3_1 _06594_ (.A(net236),
    .B(net243),
    .C(net244),
    .X(_03886_));
 sky130_fd_sc_hd__nand2_2 _06595_ (.A(_02503_),
    .B(_03886_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_2 _06596_ (.A(_03875_),
    .B(_03897_),
    .Y(_03908_));
 sky130_fd_sc_hd__xor2_4 _06597_ (.A(_03842_),
    .B(_03908_),
    .X(_03919_));
 sky130_fd_sc_hd__xnor2_1 _06598_ (.A(_02525_),
    .B(_03919_),
    .Y(_03930_));
 sky130_fd_sc_hd__clkbuf_4 _06599_ (.A(net200),
    .X(_03941_));
 sky130_fd_sc_hd__and2_2 _06600_ (.A(_03941_),
    .B(_02448_),
    .X(_03952_));
 sky130_fd_sc_hd__nor2_1 _06601_ (.A(_03930_),
    .B(_03952_),
    .Y(_03963_));
 sky130_fd_sc_hd__and2_1 _06602_ (.A(_03930_),
    .B(_03952_),
    .X(_03974_));
 sky130_fd_sc_hd__nor2_1 _06603_ (.A(_03963_),
    .B(_03974_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _06604_ (.A(_03776_),
    .B(_03985_),
    .Y(_03996_));
 sky130_fd_sc_hd__or2_1 _06605_ (.A(_03776_),
    .B(_03985_),
    .X(_04007_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(_03996_),
    .B(_04007_),
    .Y(_04018_));
 sky130_fd_sc_hd__or2_1 _06607_ (.A(_02602_),
    .B(_04018_),
    .X(_04029_));
 sky130_fd_sc_hd__nand2_1 _06608_ (.A(_02602_),
    .B(_04018_),
    .Y(_04040_));
 sky130_fd_sc_hd__and2_1 _06609_ (.A(_04029_),
    .B(_04040_),
    .X(_04051_));
 sky130_fd_sc_hd__nand3_1 _06610_ (.A(_03710_),
    .B(_03721_),
    .C(_04051_),
    .Y(_04062_));
 sky130_fd_sc_hd__a21o_1 _06611_ (.A1(_03710_),
    .A2(_03721_),
    .B1(_04051_),
    .X(_04073_));
 sky130_fd_sc_hd__nand3_2 _06612_ (.A(_02976_),
    .B(_04062_),
    .C(_04073_),
    .Y(_04084_));
 sky130_fd_sc_hd__a21o_1 _06613_ (.A1(_04062_),
    .A2(_04073_),
    .B1(_02976_),
    .X(_04095_));
 sky130_fd_sc_hd__buf_2 _06614_ (.A(net209),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_1 _06615_ (.A(_02459_),
    .B(_04106_),
    .Y(_04117_));
 sky130_fd_sc_hd__buf_2 _06616_ (.A(net140),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_4 _06617_ (.A(net149),
    .X(_04139_));
 sky130_fd_sc_hd__and3_1 _06618_ (.A(_04128_),
    .B(_02383_),
    .C(_04139_),
    .X(_04150_));
 sky130_fd_sc_hd__a22o_1 _06619_ (.A1(_04128_),
    .A2(_02383_),
    .B1(_04139_),
    .B2(_02394_),
    .X(_04161_));
 sky130_fd_sc_hd__a21bo_1 _06620_ (.A1(_02394_),
    .A2(_04150_),
    .B1_N(_04161_),
    .X(_04172_));
 sky130_fd_sc_hd__or2_1 _06621_ (.A(_04117_),
    .B(_04172_),
    .X(_04183_));
 sky130_fd_sc_hd__nand2_1 _06622_ (.A(_04117_),
    .B(_04172_),
    .Y(_04194_));
 sky130_fd_sc_hd__and2_2 _06623_ (.A(_04183_),
    .B(_04194_),
    .X(_04205_));
 sky130_fd_sc_hd__xor2_1 _06624_ (.A(_02536_),
    .B(_04205_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_2 _06625_ (.A(net158),
    .X(_04227_));
 sky130_fd_sc_hd__buf_2 _06626_ (.A(net166),
    .X(_04238_));
 sky130_fd_sc_hd__a22oi_1 _06627_ (.A1(_04227_),
    .A2(_02317_),
    .B1(_04238_),
    .B2(_02328_),
    .Y(_04249_));
 sky130_fd_sc_hd__and3_1 _06628_ (.A(_04227_),
    .B(_02317_),
    .C(_04238_),
    .X(_04259_));
 sky130_fd_sc_hd__and2_1 _06629_ (.A(_02328_),
    .B(_04259_),
    .X(_04270_));
 sky130_fd_sc_hd__or2_1 _06630_ (.A(_04249_),
    .B(_04270_),
    .X(_04281_));
 sky130_fd_sc_hd__buf_4 _06631_ (.A(net86),
    .X(_04292_));
 sky130_fd_sc_hd__buf_2 _06632_ (.A(net122),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_4 _06633_ (.A(net131),
    .X(_04314_));
 sky130_fd_sc_hd__a22o_2 _06634_ (.A1(_04303_),
    .A2(_02218_),
    .B1(_04314_),
    .B2(_02229_),
    .X(_04325_));
 sky130_fd_sc_hd__and3_2 _06635_ (.A(_04303_),
    .B(_02218_),
    .C(_04314_),
    .X(_04336_));
 sky130_fd_sc_hd__nand2_4 _06636_ (.A(_02229_),
    .B(_04336_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand4_4 _06637_ (.A(_04292_),
    .B(_02240_),
    .C(_04325_),
    .D(_04347_),
    .Y(_04358_));
 sky130_fd_sc_hd__a22o_1 _06638_ (.A1(_04292_),
    .A2(_02240_),
    .B1(_04325_),
    .B2(_04347_),
    .X(_04369_));
 sky130_fd_sc_hd__and3_1 _06639_ (.A(_02273_),
    .B(_04358_),
    .C(_04369_),
    .X(_04380_));
 sky130_fd_sc_hd__inv_2 _06640_ (.A(_04380_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21o_1 _06641_ (.A1(_04358_),
    .A2(_04369_),
    .B1(_02273_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_4 _06642_ (.A(net95),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_4 _06643_ (.A(_04413_),
    .X(_04424_));
 sky130_fd_sc_hd__buf_2 _06644_ (.A(net16),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_4 _06645_ (.A(net25),
    .X(_04446_));
 sky130_fd_sc_hd__a22o_1 _06646_ (.A1(_04435_),
    .A2(_02196_),
    .B1(_04446_),
    .B2(_02207_),
    .X(_04457_));
 sky130_fd_sc_hd__and3_1 _06647_ (.A(_04435_),
    .B(_02196_),
    .C(_04446_),
    .X(_04468_));
 sky130_fd_sc_hd__nand2_1 _06648_ (.A(_02207_),
    .B(_04468_),
    .Y(_04479_));
 sky130_fd_sc_hd__and4_1 _06649_ (.A(_02251_),
    .B(_04424_),
    .C(_04457_),
    .D(_04479_),
    .X(_04490_));
 sky130_fd_sc_hd__a22oi_1 _06650_ (.A1(_02251_),
    .A2(_04424_),
    .B1(_04457_),
    .B2(_04479_),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_1 _06651_ (.A(_04490_),
    .B(_04501_),
    .Y(_04512_));
 sky130_fd_sc_hd__and3_1 _06652_ (.A(_04391_),
    .B(_04402_),
    .C(_04512_),
    .X(_04523_));
 sky130_fd_sc_hd__a21oi_1 _06653_ (.A1(_04391_),
    .A2(_04402_),
    .B1(_04512_),
    .Y(_04534_));
 sky130_fd_sc_hd__or2_1 _06654_ (.A(_04523_),
    .B(_04534_),
    .X(_04545_));
 sky130_fd_sc_hd__nor2_1 _06655_ (.A(_02295_),
    .B(_04545_),
    .Y(_04556_));
 sky130_fd_sc_hd__and2_1 _06656_ (.A(_02295_),
    .B(_04545_),
    .X(_04567_));
 sky130_fd_sc_hd__or2_1 _06657_ (.A(_04556_),
    .B(_04567_),
    .X(_04578_));
 sky130_fd_sc_hd__xor2_1 _06658_ (.A(_04281_),
    .B(_04578_),
    .X(_04589_));
 sky130_fd_sc_hd__xnor2_1 _06659_ (.A(_04216_),
    .B(_04589_),
    .Y(_04600_));
 sky130_fd_sc_hd__xnor2_1 _06660_ (.A(_02415_),
    .B(_04600_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand3_2 _06661_ (.A(_04084_),
    .B(_04095_),
    .C(_04611_),
    .Y(_04622_));
 sky130_fd_sc_hd__a21o_1 _06662_ (.A1(_04084_),
    .A2(_04095_),
    .B1(_04611_),
    .X(_04633_));
 sky130_fd_sc_hd__nand2_1 _06663_ (.A(_04622_),
    .B(_04633_),
    .Y(_04644_));
 sky130_fd_sc_hd__xnor2_2 _06664_ (.A(_03073_),
    .B(_04644_),
    .Y(_04655_));
 sky130_fd_sc_hd__xor2_2 _06665_ (.A(_02350_),
    .B(_04655_),
    .X(_04666_));
 sky130_fd_sc_hd__xnor2_1 _06666_ (.A(net269),
    .B(_04666_),
    .Y(_04677_));
 sky130_fd_sc_hd__or2_1 _06667_ (.A(_03042_),
    .B(_04677_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_1 _06668_ (.A(_03042_),
    .B(_04677_),
    .Y(_04699_));
 sky130_fd_sc_hd__and3_1 _06669_ (.A(_02185_),
    .B(_04688_),
    .C(_04699_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _06670_ (.A(_04710_),
    .X(_00001_));
 sky130_fd_sc_hd__nand3_2 _06671_ (.A(_03216_),
    .B(_03249_),
    .C(_03271_),
    .Y(_04730_));
 sky130_fd_sc_hd__buf_2 _06672_ (.A(net228),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_4 _06673_ (.A(net219),
    .X(_04752_));
 sky130_fd_sc_hd__a22o_1 _06674_ (.A1(_03227_),
    .A2(_03260_),
    .B1(_04752_),
    .B2(_02855_),
    .X(_04763_));
 sky130_fd_sc_hd__and2_1 _06675_ (.A(net217),
    .B(_03238_),
    .X(_04774_));
 sky130_fd_sc_hd__nand2_2 _06676_ (.A(_04752_),
    .B(_03238_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_1 _06677_ (.A(_04774_),
    .B(_04785_),
    .Y(_04796_));
 sky130_fd_sc_hd__and2_1 _06678_ (.A(_04763_),
    .B(_04796_),
    .X(_04807_));
 sky130_fd_sc_hd__and3_1 _06679_ (.A(_02866_),
    .B(_04741_),
    .C(_04807_),
    .X(_04818_));
 sky130_fd_sc_hd__o21a_1 _06680_ (.A1(_04774_),
    .A2(_04785_),
    .B1(_04807_),
    .X(_04829_));
 sky130_fd_sc_hd__a21oi_1 _06681_ (.A1(_02866_),
    .A2(_04741_),
    .B1(_04829_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _06682_ (.A(_04818_),
    .B(_04840_),
    .Y(_04851_));
 sky130_fd_sc_hd__clkbuf_4 _06683_ (.A(net43),
    .X(_04862_));
 sky130_fd_sc_hd__a22oi_2 _06684_ (.A1(_03084_),
    .A2(_03194_),
    .B1(_04862_),
    .B2(_02822_),
    .Y(_04873_));
 sky130_fd_sc_hd__and4_1 _06685_ (.A(_03084_),
    .B(_02822_),
    .C(_03194_),
    .D(_04862_),
    .X(_04884_));
 sky130_fd_sc_hd__nor2_2 _06686_ (.A(_04873_),
    .B(_04884_),
    .Y(_04895_));
 sky130_fd_sc_hd__clkbuf_4 _06687_ (.A(net35),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_2 _06688_ (.A(_02811_),
    .B(_04906_),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_2 _06689_ (.A(net1),
    .B(net12),
    .Y(_04928_));
 sky130_fd_sc_hd__buf_2 _06690_ (.A(net179),
    .X(_04939_));
 sky130_fd_sc_hd__a22o_1 _06691_ (.A1(net112),
    .A2(net256),
    .B1(net179),
    .B2(net245),
    .X(_04950_));
 sky130_fd_sc_hd__a21bo_1 _06692_ (.A1(_04939_),
    .A2(_03128_),
    .B1_N(_04950_),
    .X(_04961_));
 sky130_fd_sc_hd__xor2_4 _06693_ (.A(_04928_),
    .B(_04961_),
    .X(_04972_));
 sky130_fd_sc_hd__xnor2_4 _06694_ (.A(_03139_),
    .B(_04972_),
    .Y(_04983_));
 sky130_fd_sc_hd__xnor2_4 _06695_ (.A(_04917_),
    .B(_04983_),
    .Y(_04994_));
 sky130_fd_sc_hd__xor2_4 _06696_ (.A(_03150_),
    .B(_04994_),
    .X(_05005_));
 sky130_fd_sc_hd__xnor2_4 _06697_ (.A(_04895_),
    .B(_05005_),
    .Y(_05016_));
 sky130_fd_sc_hd__and2_1 _06698_ (.A(_02844_),
    .B(_03172_),
    .X(_05027_));
 sky130_fd_sc_hd__a31o_2 _06699_ (.A1(_02822_),
    .A2(_03194_),
    .A3(_03183_),
    .B1(_05027_),
    .X(_05038_));
 sky130_fd_sc_hd__xnor2_2 _06700_ (.A(_05016_),
    .B(_05038_),
    .Y(_05049_));
 sky130_fd_sc_hd__xor2_2 _06701_ (.A(_04851_),
    .B(_05049_),
    .X(_05060_));
 sky130_fd_sc_hd__xor2_1 _06702_ (.A(_04730_),
    .B(_05060_),
    .X(_05071_));
 sky130_fd_sc_hd__and4_1 _06703_ (.A(_03337_),
    .B(_02712_),
    .C(_03348_),
    .D(_02723_),
    .X(_05082_));
 sky130_fd_sc_hd__buf_2 _06704_ (.A(net193),
    .X(_05093_));
 sky130_fd_sc_hd__a22o_1 _06705_ (.A1(net183),
    .A2(_03348_),
    .B1(net184),
    .B2(_02712_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_4 _06706_ (.A(net184),
    .X(_05115_));
 sky130_fd_sc_hd__nand4_4 _06707_ (.A(_03337_),
    .B(_02712_),
    .C(_03348_),
    .D(_05115_),
    .Y(_05126_));
 sky130_fd_sc_hd__a22o_1 _06708_ (.A1(_02723_),
    .A2(_05093_),
    .B1(_05104_),
    .B2(_05126_),
    .X(_05137_));
 sky130_fd_sc_hd__nand4_2 _06709_ (.A(_02723_),
    .B(_05093_),
    .C(_05104_),
    .D(_05126_),
    .Y(_05147_));
 sky130_fd_sc_hd__and3_1 _06710_ (.A(_05082_),
    .B(_05137_),
    .C(_05147_),
    .X(_05158_));
 sky130_fd_sc_hd__a21oi_1 _06711_ (.A1(_05137_),
    .A2(_05147_),
    .B1(_05082_),
    .Y(_05169_));
 sky130_fd_sc_hd__or2_1 _06712_ (.A(_05158_),
    .B(_05169_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_4 _06713_ (.A(net100),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_4 _06714_ (.A(net175),
    .X(_05202_));
 sky130_fd_sc_hd__a22o_1 _06715_ (.A1(_03381_),
    .A2(_03392_),
    .B1(_02745_),
    .B2(_05202_),
    .X(_05213_));
 sky130_fd_sc_hd__and4_1 _06716_ (.A(net89),
    .B(_03392_),
    .C(net78),
    .D(_05202_),
    .X(_05224_));
 sky130_fd_sc_hd__inv_2 _06717_ (.A(_05224_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand4_2 _06718_ (.A(_02734_),
    .B(_05191_),
    .C(_05213_),
    .D(_05235_),
    .Y(_05246_));
 sky130_fd_sc_hd__a22o_1 _06719_ (.A1(_02734_),
    .A2(_05191_),
    .B1(_05213_),
    .B2(_05235_),
    .X(_05257_));
 sky130_fd_sc_hd__nand2_1 _06720_ (.A(_05246_),
    .B(_05257_),
    .Y(_05268_));
 sky130_fd_sc_hd__xor2_1 _06721_ (.A(_05180_),
    .B(_05268_),
    .X(_05279_));
 sky130_fd_sc_hd__and2_1 _06722_ (.A(_03436_),
    .B(_05279_),
    .X(_05290_));
 sky130_fd_sc_hd__nor2_1 _06723_ (.A(_03436_),
    .B(_05279_),
    .Y(_05301_));
 sky130_fd_sc_hd__or2_1 _06724_ (.A(_05290_),
    .B(_05301_),
    .X(_05312_));
 sky130_fd_sc_hd__or2_1 _06725_ (.A(_05071_),
    .B(_05312_),
    .X(_05323_));
 sky130_fd_sc_hd__nand2_1 _06726_ (.A(_05071_),
    .B(_05312_),
    .Y(_05334_));
 sky130_fd_sc_hd__o21ai_1 _06727_ (.A1(_03326_),
    .A2(_03491_),
    .B1(_03304_),
    .Y(_05345_));
 sky130_fd_sc_hd__and3_1 _06728_ (.A(_05323_),
    .B(_05334_),
    .C(_05345_),
    .X(_05356_));
 sky130_fd_sc_hd__a21oi_1 _06729_ (.A1(_05323_),
    .A2(_05334_),
    .B1(_05345_),
    .Y(_05367_));
 sky130_fd_sc_hd__or2_1 _06730_ (.A(_03568_),
    .B(_03634_),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_4 _06731_ (.A(net105),
    .X(_05389_));
 sky130_fd_sc_hd__a22oi_1 _06732_ (.A1(_03524_),
    .A2(_03546_),
    .B1(_05389_),
    .B2(_02635_),
    .Y(_05400_));
 sky130_fd_sc_hd__and4_1 _06733_ (.A(net104),
    .B(net113),
    .C(net114),
    .D(_05389_),
    .X(_05411_));
 sky130_fd_sc_hd__or2_1 _06734_ (.A(_05400_),
    .B(_05411_),
    .X(_05422_));
 sky130_fd_sc_hd__xnor2_1 _06735_ (.A(_03425_),
    .B(_05422_),
    .Y(_05433_));
 sky130_fd_sc_hd__clkbuf_4 _06736_ (.A(net115),
    .X(_05444_));
 sky130_fd_sc_hd__nand3_1 _06737_ (.A(net103),
    .B(_05444_),
    .C(_03535_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21a_1 _06738_ (.A1(_05444_),
    .A2(_03535_),
    .B1(_02646_),
    .X(_05466_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(_05455_),
    .B(_05466_),
    .Y(_05477_));
 sky130_fd_sc_hd__and4_1 _06740_ (.A(net69),
    .B(net76),
    .C(net77),
    .D(net70),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_4 _06741_ (.A(net70),
    .X(_05498_));
 sky130_fd_sc_hd__a22o_1 _06742_ (.A1(_03579_),
    .A2(_03590_),
    .B1(_05498_),
    .B2(_02657_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_4 _06743_ (.A(net79),
    .X(_05520_));
 sky130_fd_sc_hd__and4b_1 _06744_ (.A_N(_05487_),
    .B(_05509_),
    .C(net68),
    .D(_05520_),
    .X(_05531_));
 sky130_fd_sc_hd__inv_2 _06745_ (.A(_05487_),
    .Y(_05542_));
 sky130_fd_sc_hd__a22oi_1 _06746_ (.A1(net68),
    .A2(_05520_),
    .B1(_05542_),
    .B2(_05509_),
    .Y(_05553_));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(_05531_),
    .B(_05553_),
    .Y(_05564_));
 sky130_fd_sc_hd__xnor2_1 _06748_ (.A(_05477_),
    .B(_05564_),
    .Y(_05575_));
 sky130_fd_sc_hd__xor2_1 _06749_ (.A(_03623_),
    .B(_05575_),
    .X(_05586_));
 sky130_fd_sc_hd__or2_1 _06750_ (.A(_05433_),
    .B(_05586_),
    .X(_05597_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(_05433_),
    .B(_05586_),
    .Y(_05608_));
 sky130_fd_sc_hd__and3_1 _06752_ (.A(_03469_),
    .B(_05597_),
    .C(_05608_),
    .X(_05619_));
 sky130_fd_sc_hd__and2_1 _06753_ (.A(_05597_),
    .B(_05608_),
    .X(_05630_));
 sky130_fd_sc_hd__nor2_1 _06754_ (.A(_03469_),
    .B(_05630_),
    .Y(_05641_));
 sky130_fd_sc_hd__or2_1 _06755_ (.A(_05619_),
    .B(_05641_),
    .X(_05652_));
 sky130_fd_sc_hd__nor2_1 _06756_ (.A(_05378_),
    .B(_05652_),
    .Y(_05663_));
 sky130_fd_sc_hd__and2_1 _06757_ (.A(_05378_),
    .B(_05652_),
    .X(_05674_));
 sky130_fd_sc_hd__or2_1 _06758_ (.A(_05663_),
    .B(_05674_),
    .X(_05685_));
 sky130_fd_sc_hd__or3_2 _06759_ (.A(_05356_),
    .B(_05367_),
    .C(_05685_),
    .X(_05696_));
 sky130_fd_sc_hd__o21ai_1 _06760_ (.A1(_05356_),
    .A2(_05367_),
    .B1(_05685_),
    .Y(_05707_));
 sky130_fd_sc_hd__a21bo_1 _06761_ (.A1(_02899_),
    .A2(_03502_),
    .B1_N(_03689_),
    .X(_05718_));
 sky130_fd_sc_hd__and3_1 _06762_ (.A(_05696_),
    .B(_05707_),
    .C(_05718_),
    .X(_05729_));
 sky130_fd_sc_hd__a21oi_1 _06763_ (.A1(_05696_),
    .A2(_05707_),
    .B1(_05718_),
    .Y(_05740_));
 sky130_fd_sc_hd__clkbuf_4 _06764_ (.A(net52),
    .X(_05750_));
 sky130_fd_sc_hd__buf_2 _06765_ (.A(net61),
    .X(_05761_));
 sky130_fd_sc_hd__a22o_1 _06766_ (.A1(_03732_),
    .A2(_03743_),
    .B1(_02580_),
    .B2(_05761_),
    .X(_05772_));
 sky130_fd_sc_hd__and4_1 _06767_ (.A(_03732_),
    .B(_03743_),
    .C(_02580_),
    .D(_05761_),
    .X(_05783_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(_05783_),
    .Y(_05794_));
 sky130_fd_sc_hd__and4_1 _06769_ (.A(_02569_),
    .B(_05750_),
    .C(_05772_),
    .D(_05794_),
    .X(_05805_));
 sky130_fd_sc_hd__a22oi_1 _06770_ (.A1(_02569_),
    .A2(_05750_),
    .B1(_05772_),
    .B2(_05794_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _06771_ (.A(_05805_),
    .B(_05816_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_03765_),
    .B(_05827_),
    .Y(_05838_));
 sky130_fd_sc_hd__or2_1 _06773_ (.A(_03765_),
    .B(_05827_),
    .X(_05849_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(_05838_),
    .B(_05849_),
    .Y(_05860_));
 sky130_fd_sc_hd__or2_1 _06775_ (.A(_03842_),
    .B(_03908_),
    .X(_05871_));
 sky130_fd_sc_hd__clkbuf_4 _06776_ (.A(net8),
    .X(_05882_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(_02481_),
    .B(_05882_),
    .Y(_05893_));
 sky130_fd_sc_hd__and3b_1 _06778_ (.A_N(net252),
    .B(net254),
    .C(_03787_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_2 _06779_ (.A(net254),
    .X(_05914_));
 sky130_fd_sc_hd__a22oi_1 _06780_ (.A1(_03820_),
    .A2(_03798_),
    .B1(_05914_),
    .B2(_02470_),
    .Y(_05925_));
 sky130_fd_sc_hd__and3b_1 _06781_ (.A_N(_05914_),
    .B(_03787_),
    .C(net252),
    .X(_05936_));
 sky130_fd_sc_hd__or3_2 _06782_ (.A(_05904_),
    .B(_05925_),
    .C(_05936_),
    .X(_05947_));
 sky130_fd_sc_hd__xor2_2 _06783_ (.A(_05893_),
    .B(_05947_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_4 _06784_ (.A(net246),
    .X(_05969_));
 sky130_fd_sc_hd__buf_4 _06785_ (.A(net237),
    .X(_05980_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(_05980_),
    .B(_03886_),
    .Y(_05991_));
 sky130_fd_sc_hd__a22o_1 _06787_ (.A1(_03853_),
    .A2(_03864_),
    .B1(_05980_),
    .B2(_02492_),
    .X(_06001_));
 sky130_fd_sc_hd__and4_1 _06788_ (.A(net235),
    .B(_05969_),
    .C(_05991_),
    .D(_06001_),
    .X(_06012_));
 sky130_fd_sc_hd__a22oi_1 _06789_ (.A1(_02503_),
    .A2(_05969_),
    .B1(_05991_),
    .B2(_06001_),
    .Y(_06023_));
 sky130_fd_sc_hd__nor2_1 _06790_ (.A(_06012_),
    .B(_06023_),
    .Y(_06034_));
 sky130_fd_sc_hd__xnor2_2 _06791_ (.A(_03897_),
    .B(_06034_),
    .Y(_06045_));
 sky130_fd_sc_hd__xnor2_2 _06792_ (.A(_05958_),
    .B(_06045_),
    .Y(_06055_));
 sky130_fd_sc_hd__xor2_2 _06793_ (.A(_05871_),
    .B(_06055_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_4 _06794_ (.A(net202),
    .X(_06077_));
 sky130_fd_sc_hd__clkbuf_4 _06795_ (.A(_06077_),
    .X(_06086_));
 sky130_fd_sc_hd__nand2_1 _06796_ (.A(_02448_),
    .B(_06086_),
    .Y(_06095_));
 sky130_fd_sc_hd__xor2_2 _06797_ (.A(_06066_),
    .B(_06095_),
    .X(_06104_));
 sky130_fd_sc_hd__nor2_1 _06798_ (.A(_05860_),
    .B(_06104_),
    .Y(_06112_));
 sky130_fd_sc_hd__and2_1 _06799_ (.A(_05860_),
    .B(_06104_),
    .X(_06114_));
 sky130_fd_sc_hd__nor2_1 _06800_ (.A(_06112_),
    .B(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__and2_1 _06801_ (.A(_03656_),
    .B(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__nor2_1 _06802_ (.A(_03656_),
    .B(_06115_),
    .Y(_06117_));
 sky130_fd_sc_hd__or2_1 _06803_ (.A(_06116_),
    .B(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__nor2_1 _06804_ (.A(_03996_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__and2_1 _06805_ (.A(_03996_),
    .B(_06118_),
    .X(_06120_));
 sky130_fd_sc_hd__or2_1 _06806_ (.A(_06119_),
    .B(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__or3_2 _06807_ (.A(_05729_),
    .B(_05740_),
    .C(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__o21ai_1 _06808_ (.A1(_05729_),
    .A2(_05740_),
    .B1(_06121_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _06809_ (.A(_03710_),
    .B(_04062_),
    .Y(_06124_));
 sky130_fd_sc_hd__and3_1 _06810_ (.A(_06122_),
    .B(_06123_),
    .C(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__a21oi_1 _06811_ (.A1(_06122_),
    .A2(_06123_),
    .B1(_06124_),
    .Y(_06126_));
 sky130_fd_sc_hd__buf_2 _06812_ (.A(net159),
    .X(_06127_));
 sky130_fd_sc_hd__a22o_1 _06813_ (.A1(_04227_),
    .A2(_04238_),
    .B1(_06127_),
    .B2(_02317_),
    .X(_06128_));
 sky130_fd_sc_hd__a21bo_1 _06814_ (.A1(_06127_),
    .A2(_04259_),
    .B1_N(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_4 _06815_ (.A(net168),
    .X(_06130_));
 sky130_fd_sc_hd__nand2_1 _06816_ (.A(_02328_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__xor2_2 _06817_ (.A(_06129_),
    .B(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__xnor2_1 _06818_ (.A(_04490_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__clkbuf_4 _06819_ (.A(net96),
    .X(_06134_));
 sky130_fd_sc_hd__a22oi_1 _06820_ (.A1(_04292_),
    .A2(_04424_),
    .B1(_06134_),
    .B2(_02251_),
    .Y(_06135_));
 sky130_fd_sc_hd__and4_1 _06821_ (.A(_04292_),
    .B(_02251_),
    .C(_04424_),
    .D(_06134_),
    .X(_06136_));
 sky130_fd_sc_hd__nor2_1 _06822_ (.A(_06135_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__clkbuf_4 _06823_ (.A(net17),
    .X(_06138_));
 sky130_fd_sc_hd__a22oi_1 _06824_ (.A1(_04435_),
    .A2(_04446_),
    .B1(_06138_),
    .B2(_02196_),
    .Y(_06139_));
 sky130_fd_sc_hd__and2_1 _06825_ (.A(_06138_),
    .B(_04468_),
    .X(_06140_));
 sky130_fd_sc_hd__or2_1 _06826_ (.A(_06139_),
    .B(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_4 _06827_ (.A(net26),
    .X(_06142_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(_02207_),
    .B(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__mux2_1 _06829_ (.A0(_06142_),
    .A1(_06143_),
    .S(_04479_),
    .X(_06144_));
 sky130_fd_sc_hd__nor2_1 _06830_ (.A(_06141_),
    .B(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__and2_1 _06831_ (.A(_06141_),
    .B(_06144_),
    .X(_06146_));
 sky130_fd_sc_hd__nor2_1 _06832_ (.A(_06145_),
    .B(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__nand2_1 _06833_ (.A(_06137_),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__or2_1 _06834_ (.A(_06137_),
    .B(_06147_),
    .X(_06149_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_06148_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__buf_2 _06836_ (.A(net132),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_4 _06837_ (.A(net124),
    .X(_06152_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_06152_),
    .B(_04336_),
    .Y(_06153_));
 sky130_fd_sc_hd__a22o_1 _06839_ (.A1(_04303_),
    .A2(_04314_),
    .B1(_06152_),
    .B2(_02218_),
    .X(_06154_));
 sky130_fd_sc_hd__and4_1 _06840_ (.A(net121),
    .B(_06151_),
    .C(_06153_),
    .D(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__a22oi_1 _06841_ (.A1(_02229_),
    .A2(_06151_),
    .B1(_06153_),
    .B2(_06154_),
    .Y(_06156_));
 sky130_fd_sc_hd__nor2_2 _06842_ (.A(_06155_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__xnor2_4 _06843_ (.A(_04347_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__clkbuf_4 _06844_ (.A(net87),
    .X(_06159_));
 sky130_fd_sc_hd__nand2_2 _06845_ (.A(_02240_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__xor2_4 _06846_ (.A(_06158_),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nand2_1 _06847_ (.A(_04358_),
    .B(_04391_),
    .Y(_06162_));
 sky130_fd_sc_hd__xnor2_1 _06848_ (.A(_06161_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__xnor2_1 _06849_ (.A(_06150_),
    .B(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__xnor2_1 _06850_ (.A(_04523_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__nor2_1 _06851_ (.A(_06133_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__inv_2 _06852_ (.A(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(_06133_),
    .B(_06165_),
    .Y(_06168_));
 sky130_fd_sc_hd__and2b_1 _06854_ (.A_N(_02536_),
    .B(_04205_),
    .X(_06169_));
 sky130_fd_sc_hd__and2b_1 _06855_ (.A_N(_02525_),
    .B(_03919_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_4 _06856_ (.A(net150),
    .X(_06171_));
 sky130_fd_sc_hd__buf_2 _06857_ (.A(net210),
    .X(_06172_));
 sky130_fd_sc_hd__buf_2 _06858_ (.A(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__a22oi_1 _06859_ (.A1(_03941_),
    .A2(_04106_),
    .B1(_06173_),
    .B2(_02459_),
    .Y(_06174_));
 sky130_fd_sc_hd__and4_1 _06860_ (.A(_03941_),
    .B(_02459_),
    .C(_04106_),
    .D(_06173_),
    .X(_06175_));
 sky130_fd_sc_hd__nor2_1 _06861_ (.A(_06174_),
    .B(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__clkbuf_4 _06862_ (.A(net141),
    .X(_06177_));
 sky130_fd_sc_hd__buf_2 _06863_ (.A(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__nand3b_1 _06864_ (.A_N(_02394_),
    .B(_06178_),
    .C(_04150_),
    .Y(_06179_));
 sky130_fd_sc_hd__a22o_1 _06865_ (.A1(_04128_),
    .A2(_04139_),
    .B1(_06178_),
    .B2(_02383_),
    .X(_06180_));
 sky130_fd_sc_hd__nand3b_2 _06866_ (.A_N(_06178_),
    .B(_04150_),
    .C(_02394_),
    .Y(_06181_));
 sky130_fd_sc_hd__and4_1 _06867_ (.A(_06176_),
    .B(_06179_),
    .C(_06180_),
    .D(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__a31o_1 _06868_ (.A1(_06179_),
    .A2(_06180_),
    .A3(_06181_),
    .B1(_06176_),
    .X(_06183_));
 sky130_fd_sc_hd__or2b_1 _06869_ (.A(_06182_),
    .B_N(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__xor2_1 _06870_ (.A(_04183_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__and3_1 _06871_ (.A(_02394_),
    .B(_06171_),
    .C(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__a21oi_1 _06872_ (.A1(_02394_),
    .A2(_06171_),
    .B1(_06185_),
    .Y(_06187_));
 sky130_fd_sc_hd__nor2_2 _06873_ (.A(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__o21ai_2 _06874_ (.A1(_06170_),
    .A2(_03974_),
    .B1(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__or3_1 _06875_ (.A(_06170_),
    .B(_03974_),
    .C(_06188_),
    .X(_06190_));
 sky130_fd_sc_hd__and2_1 _06876_ (.A(_06189_),
    .B(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_06169_),
    .B(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__or2_1 _06878_ (.A(_06169_),
    .B(_06191_),
    .X(_06193_));
 sky130_fd_sc_hd__and2_1 _06879_ (.A(_06192_),
    .B(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__and3_1 _06880_ (.A(_06167_),
    .B(_06168_),
    .C(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__a21oi_1 _06881_ (.A1(_06167_),
    .A2(_06168_),
    .B1(_06194_),
    .Y(_06196_));
 sky130_fd_sc_hd__or3_2 _06882_ (.A(_04029_),
    .B(_06195_),
    .C(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__o21ai_2 _06883_ (.A1(_06195_),
    .A2(_06196_),
    .B1(_04029_),
    .Y(_06198_));
 sky130_fd_sc_hd__and2b_1 _06884_ (.A_N(_04216_),
    .B(_04589_),
    .X(_06199_));
 sky130_fd_sc_hd__a21oi_2 _06885_ (.A1(_06197_),
    .A2(_06198_),
    .B1(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__nand3_2 _06886_ (.A(_06199_),
    .B(_06197_),
    .C(_06198_),
    .Y(_06201_));
 sky130_fd_sc_hd__inv_2 _06887_ (.A(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor4_2 _06888_ (.A(_06125_),
    .B(_06126_),
    .C(_06200_),
    .D(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__o22a_1 _06889_ (.A1(_06125_),
    .A2(_06126_),
    .B1(_06200_),
    .B2(_06202_),
    .X(_06204_));
 sky130_fd_sc_hd__a211oi_1 _06890_ (.A1(_04084_),
    .A2(_04622_),
    .B1(_06203_),
    .C1(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__o211a_1 _06891_ (.A1(_06203_),
    .A2(_06204_),
    .B1(_04084_),
    .C1(_04622_),
    .X(_06206_));
 sky130_fd_sc_hd__or2b_1 _06892_ (.A(_02415_),
    .B_N(_04600_),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_1 _06893_ (.A(_04270_),
    .B(_04556_),
    .Y(_06208_));
 sky130_fd_sc_hd__or2_1 _06894_ (.A(_04270_),
    .B(_04556_),
    .X(_06209_));
 sky130_fd_sc_hd__a2bb2o_1 _06895_ (.A1_N(_04281_),
    .A2_N(_04578_),
    .B1(_06208_),
    .B2(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__or2b_2 _06896_ (.A(_06207_),
    .B_N(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__or2b_1 _06897_ (.A(_06210_),
    .B_N(_06207_),
    .X(_06212_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(_06211_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__or3_2 _06899_ (.A(_06205_),
    .B(_06206_),
    .C(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__o21ai_1 _06900_ (.A1(_06205_),
    .A2(_06206_),
    .B1(_06213_),
    .Y(_06215_));
 sky130_fd_sc_hd__and2_1 _06901_ (.A(_06214_),
    .B(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__a32o_1 _06902_ (.A1(_03073_),
    .A2(_04622_),
    .A3(_04633_),
    .B1(_04655_),
    .B2(_02350_),
    .X(_06217_));
 sky130_fd_sc_hd__xor2_2 _06903_ (.A(_06216_),
    .B(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__xnor2_1 _06904_ (.A(net278),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__a21boi_1 _06905_ (.A1(net269),
    .A2(_04666_),
    .B1_N(_04688_),
    .Y(_06220_));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(_06219_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__or2_1 _06907_ (.A(_06219_),
    .B(_06220_),
    .X(_06222_));
 sky130_fd_sc_hd__and3_1 _06908_ (.A(_02185_),
    .B(_06221_),
    .C(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _06909_ (.A(_06223_),
    .X(_00002_));
 sky130_fd_sc_hd__and2_1 _06910_ (.A(_06216_),
    .B(_06217_),
    .X(_06224_));
 sky130_fd_sc_hd__a211o_1 _06911_ (.A1(_04084_),
    .A2(_04622_),
    .B1(_06203_),
    .C1(_06204_),
    .X(_06225_));
 sky130_fd_sc_hd__a21o_1 _06912_ (.A1(_04523_),
    .A2(_06164_),
    .B1(_06166_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_4 _06913_ (.A(net169),
    .X(_06227_));
 sky130_fd_sc_hd__a32o_1 _06914_ (.A1(_02328_),
    .A2(_06130_),
    .A3(_06128_),
    .B1(_04259_),
    .B2(_06127_),
    .X(_06228_));
 sky130_fd_sc_hd__and3_1 _06915_ (.A(_02328_),
    .B(_06227_),
    .C(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__a21oi_1 _06916_ (.A1(_02328_),
    .A2(_06227_),
    .B1(_06228_),
    .Y(_06230_));
 sky130_fd_sc_hd__nor2_1 _06917_ (.A(_06229_),
    .B(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__and3_1 _06918_ (.A(_04490_),
    .B(_06132_),
    .C(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__a21oi_1 _06919_ (.A1(_04490_),
    .A2(_06132_),
    .B1(_06231_),
    .Y(_06233_));
 sky130_fd_sc_hd__nor2_1 _06920_ (.A(_06232_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__xnor2_1 _06921_ (.A(_06226_),
    .B(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__a21oi_2 _06922_ (.A1(_06197_),
    .A2(_06201_),
    .B1(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__and3_1 _06923_ (.A(_06197_),
    .B(_06201_),
    .C(_06235_),
    .X(_06237_));
 sky130_fd_sc_hd__or2_1 _06924_ (.A(_06236_),
    .B(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__and2_1 _06925_ (.A(_06208_),
    .B(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__nor2_2 _06926_ (.A(_06208_),
    .B(_06238_),
    .Y(_06240_));
 sky130_fd_sc_hd__nor2_1 _06927_ (.A(_06239_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__inv_2 _06928_ (.A(_06195_),
    .Y(_06242_));
 sky130_fd_sc_hd__clkbuf_4 _06929_ (.A(net160),
    .X(_06243_));
 sky130_fd_sc_hd__a22oi_2 _06930_ (.A1(_04238_),
    .A2(_06127_),
    .B1(_06243_),
    .B2(_02317_),
    .Y(_06244_));
 sky130_fd_sc_hd__and4_1 _06931_ (.A(_02317_),
    .B(_04238_),
    .C(_06127_),
    .D(_06243_),
    .X(_06245_));
 sky130_fd_sc_hd__nand2_1 _06932_ (.A(_04227_),
    .B(_06130_),
    .Y(_06246_));
 sky130_fd_sc_hd__o21a_1 _06933_ (.A1(_06244_),
    .A2(_06245_),
    .B1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__nor3_1 _06934_ (.A(_06244_),
    .B(_06245_),
    .C(_06246_),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _06935_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__a31o_1 _06936_ (.A1(_02207_),
    .A2(_06142_),
    .A3(_04468_),
    .B1(_06145_),
    .X(_06250_));
 sky130_fd_sc_hd__xnor2_2 _06937_ (.A(_06249_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__xor2_1 _06938_ (.A(_06148_),
    .B(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__buf_2 _06939_ (.A(net97),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_4 _06940_ (.A(net96),
    .X(_06254_));
 sky130_fd_sc_hd__nand4_1 _06941_ (.A(net86),
    .B(_04413_),
    .C(net87),
    .D(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__a22o_1 _06942_ (.A1(_04413_),
    .A2(net87),
    .B1(_06254_),
    .B2(net86),
    .X(_06256_));
 sky130_fd_sc_hd__and4_1 _06943_ (.A(net85),
    .B(_06253_),
    .C(_06255_),
    .D(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__a22oi_1 _06944_ (.A1(_02251_),
    .A2(_06253_),
    .B1(_06255_),
    .B2(_06256_),
    .Y(_06258_));
 sky130_fd_sc_hd__nor2_1 _06945_ (.A(_06257_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_1 _06946_ (.A(_06136_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__clkbuf_4 _06947_ (.A(net18),
    .X(_06261_));
 sky130_fd_sc_hd__a22oi_2 _06948_ (.A1(_04446_),
    .A2(_06138_),
    .B1(_06261_),
    .B2(_02196_),
    .Y(_06262_));
 sky130_fd_sc_hd__and4_1 _06949_ (.A(net24),
    .B(net25),
    .C(_06138_),
    .D(_06261_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_4 _06950_ (.A(net27),
    .X(_06264_));
 sky130_fd_sc_hd__nand4_2 _06951_ (.A(_04435_),
    .B(_02207_),
    .C(_06142_),
    .D(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__a22o_1 _06952_ (.A1(_04435_),
    .A2(_06142_),
    .B1(_06264_),
    .B2(_02207_),
    .X(_06266_));
 sky130_fd_sc_hd__and3_1 _06953_ (.A(_06140_),
    .B(_06265_),
    .C(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__a21oi_1 _06954_ (.A1(_06265_),
    .A2(_06266_),
    .B1(_06140_),
    .Y(_06268_));
 sky130_fd_sc_hd__nor4_1 _06955_ (.A(_06262_),
    .B(_06263_),
    .C(_06267_),
    .D(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__o22a_1 _06956_ (.A1(_06262_),
    .A2(_06263_),
    .B1(_06267_),
    .B2(_06268_),
    .X(_06270_));
 sky130_fd_sc_hd__nor2_1 _06957_ (.A(net308),
    .B(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__xnor2_1 _06958_ (.A(_06260_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__and3_2 _06959_ (.A(_02229_),
    .B(_04336_),
    .C(_06157_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_2 _06960_ (.A(net125),
    .X(_06274_));
 sky130_fd_sc_hd__nand4_1 _06961_ (.A(_02218_),
    .B(_04314_),
    .C(_06152_),
    .D(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__a22o_1 _06962_ (.A1(_04314_),
    .A2(net124),
    .B1(net125),
    .B2(_02218_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_2 _06963_ (.A(_06275_),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__and2_2 _06964_ (.A(_04303_),
    .B(net132),
    .X(_06278_));
 sky130_fd_sc_hd__xor2_4 _06965_ (.A(_06277_),
    .B(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a32o_2 _06966_ (.A1(net121),
    .A2(_06151_),
    .A3(_06154_),
    .B1(_04336_),
    .B2(_06152_),
    .X(_06280_));
 sky130_fd_sc_hd__xor2_4 _06967_ (.A(_06279_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__xor2_4 _06968_ (.A(_06273_),
    .B(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_4 _06969_ (.A(net133),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_4 _06970_ (.A(net88),
    .X(_06284_));
 sky130_fd_sc_hd__a22o_1 _06971_ (.A1(_02229_),
    .A2(_06283_),
    .B1(_06284_),
    .B2(_02240_),
    .X(_06285_));
 sky130_fd_sc_hd__nand4_4 _06972_ (.A(_02229_),
    .B(_02240_),
    .C(_06283_),
    .D(_06284_),
    .Y(_06286_));
 sky130_fd_sc_hd__and2_2 _06973_ (.A(_06285_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__xnor2_4 _06974_ (.A(_06282_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__nand3_2 _06975_ (.A(_02240_),
    .B(_06159_),
    .C(_06158_),
    .Y(_06289_));
 sky130_fd_sc_hd__o21a_1 _06976_ (.A1(_04358_),
    .A2(_06161_),
    .B1(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__xnor2_1 _06977_ (.A(_06288_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(_06272_),
    .B(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__or2_1 _06979_ (.A(_06272_),
    .B(_06291_),
    .X(_06293_));
 sky130_fd_sc_hd__nand2_1 _06980_ (.A(_06292_),
    .B(_06293_),
    .Y(_06294_));
 sky130_fd_sc_hd__or2b_1 _06981_ (.A(_06150_),
    .B_N(_06163_),
    .X(_06295_));
 sky130_fd_sc_hd__o21a_1 _06982_ (.A1(_04391_),
    .A2(_06161_),
    .B1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__or2_1 _06983_ (.A(_06294_),
    .B(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__nand2_1 _06984_ (.A(_06294_),
    .B(_06296_),
    .Y(_06298_));
 sky130_fd_sc_hd__and3_1 _06985_ (.A(_06252_),
    .B(_06297_),
    .C(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__a21oi_1 _06986_ (.A1(_06297_),
    .A2(_06298_),
    .B1(_06252_),
    .Y(_06300_));
 sky130_fd_sc_hd__nor2_1 _06987_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__nor2_1 _06988_ (.A(_05871_),
    .B(_06055_),
    .Y(_06302_));
 sky130_fd_sc_hd__and3_1 _06989_ (.A(_02448_),
    .B(_06086_),
    .C(_06066_),
    .X(_06303_));
 sky130_fd_sc_hd__buf_2 _06990_ (.A(net211),
    .X(_06304_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(_02459_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__and3_1 _06992_ (.A(net200),
    .B(net209),
    .C(_06172_),
    .X(_06306_));
 sky130_fd_sc_hd__a22o_1 _06993_ (.A1(net209),
    .A2(net202),
    .B1(_06172_),
    .B2(net200),
    .X(_06307_));
 sky130_fd_sc_hd__a21bo_1 _06994_ (.A1(_06086_),
    .A2(_06306_),
    .B1_N(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__xor2_1 _06995_ (.A(_06305_),
    .B(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__xnor2_1 _06996_ (.A(_06175_),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__clkbuf_4 _06997_ (.A(net142),
    .X(_06311_));
 sky130_fd_sc_hd__nand4_2 _06998_ (.A(_02383_),
    .B(_04139_),
    .C(_06177_),
    .D(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__a21o_1 _06999_ (.A1(_06178_),
    .A2(_04150_),
    .B1(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__a22o_1 _07000_ (.A1(_04139_),
    .A2(_06178_),
    .B1(_06311_),
    .B2(_02383_),
    .X(_06314_));
 sky130_fd_sc_hd__nand3_1 _07001_ (.A(_06178_),
    .B(_04150_),
    .C(_06312_),
    .Y(_06315_));
 sky130_fd_sc_hd__nand3_1 _07002_ (.A(_06313_),
    .B(_06314_),
    .C(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__xor2_1 _07003_ (.A(_06310_),
    .B(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__xnor2_1 _07004_ (.A(_06182_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__clkbuf_4 _07005_ (.A(net151),
    .X(_06319_));
 sky130_fd_sc_hd__a22o_1 _07006_ (.A1(_04128_),
    .A2(_06171_),
    .B1(_06319_),
    .B2(_02394_),
    .X(_06320_));
 sky130_fd_sc_hd__inv_2 _07007_ (.A(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__and4_1 _07008_ (.A(_04128_),
    .B(net139),
    .C(_06171_),
    .D(_06319_),
    .X(_06322_));
 sky130_fd_sc_hd__nor3_2 _07009_ (.A(_06181_),
    .B(_06321_),
    .C(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__o21a_1 _07010_ (.A1(_06321_),
    .A2(_06322_),
    .B1(_06181_),
    .X(_06324_));
 sky130_fd_sc_hd__or2_1 _07011_ (.A(_06323_),
    .B(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__or2_1 _07012_ (.A(_06318_),
    .B(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__nand2_1 _07013_ (.A(_06318_),
    .B(_06325_),
    .Y(_06327_));
 sky130_fd_sc_hd__and2_2 _07014_ (.A(_06326_),
    .B(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__o21ba_2 _07015_ (.A1(_04183_),
    .A2(_06184_),
    .B1_N(_06186_),
    .X(_06329_));
 sky130_fd_sc_hd__xnor2_4 _07016_ (.A(_06328_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ai_4 _07017_ (.A1(_06302_),
    .A2(_06303_),
    .B1(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__or3_2 _07018_ (.A(_06302_),
    .B(_06303_),
    .C(_06330_),
    .X(_06332_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_06331_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__xnor2_1 _07020_ (.A(_06189_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__inv_2 _07021_ (.A(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_1 _07022_ (.A(_06301_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__o21ba_1 _07023_ (.A1(_06116_),
    .A2(_06119_),
    .B1_N(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__nor3b_1 _07024_ (.A(_06116_),
    .B(_06119_),
    .C_N(_06336_),
    .Y(_06338_));
 sky130_fd_sc_hd__a211oi_2 _07025_ (.A1(_06192_),
    .A2(_06242_),
    .B1(_06337_),
    .C1(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__o211a_1 _07026_ (.A1(_06337_),
    .A2(_06338_),
    .B1(_06192_),
    .C1(_06242_),
    .X(_06340_));
 sky130_fd_sc_hd__inv_2 _07027_ (.A(_06122_),
    .Y(_06341_));
 sky130_fd_sc_hd__and3_1 _07028_ (.A(_02668_),
    .B(_03612_),
    .C(_05575_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_4 _07029_ (.A(net53),
    .X(_06343_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(_02569_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__and4_1 _07031_ (.A(net51),
    .B(net60),
    .C(net52),
    .D(net61),
    .X(_06345_));
 sky130_fd_sc_hd__a22o_1 _07032_ (.A1(net60),
    .A2(net52),
    .B1(net61),
    .B2(net51),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_4 _07033_ (.A(net62),
    .X(_06347_));
 sky130_fd_sc_hd__and4b_1 _07034_ (.A_N(_06345_),
    .B(_06346_),
    .C(net50),
    .D(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__inv_2 _07035_ (.A(_06345_),
    .Y(_06349_));
 sky130_fd_sc_hd__a22o_1 _07036_ (.A1(_02580_),
    .A2(_06347_),
    .B1(_06349_),
    .B2(_06346_),
    .X(_06350_));
 sky130_fd_sc_hd__and2b_1 _07037_ (.A_N(_06348_),
    .B(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__xnor2_1 _07038_ (.A(_06344_),
    .B(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__and2_1 _07039_ (.A(_05783_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nand2_1 _07040_ (.A(_05805_),
    .B(_06352_),
    .Y(_06354_));
 sky130_fd_sc_hd__or2_1 _07041_ (.A(_05805_),
    .B(_06352_),
    .X(_06355_));
 sky130_fd_sc_hd__a21oi_1 _07042_ (.A1(_06354_),
    .A2(_06355_),
    .B1(_05783_),
    .Y(_06356_));
 sky130_fd_sc_hd__or3_2 _07043_ (.A(_05838_),
    .B(_06353_),
    .C(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__o21ai_2 _07044_ (.A1(_06353_),
    .A2(_06356_),
    .B1(_05838_),
    .Y(_06358_));
 sky130_fd_sc_hd__and3_2 _07045_ (.A(_06342_),
    .B(_06357_),
    .C(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__a21oi_1 _07046_ (.A1(_06357_),
    .A2(_06358_),
    .B1(_06342_),
    .Y(_06360_));
 sky130_fd_sc_hd__buf_2 _07047_ (.A(net203),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_4 _07048_ (.A(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(_02448_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__or4_2 _07050_ (.A(_03897_),
    .B(_06012_),
    .C(_06023_),
    .D(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__a32o_1 _07051_ (.A1(_02503_),
    .A2(_03886_),
    .A3(_06034_),
    .B1(_02448_),
    .B2(_06362_),
    .X(_06365_));
 sky130_fd_sc_hd__and2_1 _07052_ (.A(_06364_),
    .B(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(_05958_),
    .B(_06045_),
    .Y(_06367_));
 sky130_fd_sc_hd__buf_4 _07054_ (.A(net9),
    .X(_06368_));
 sky130_fd_sc_hd__a22o_1 _07055_ (.A1(_03820_),
    .A2(_05882_),
    .B1(_06368_),
    .B2(net252),
    .X(_06369_));
 sky130_fd_sc_hd__and4_1 _07056_ (.A(net253),
    .B(net252),
    .C(net8),
    .D(net9),
    .X(_06370_));
 sky130_fd_sc_hd__inv_2 _07057_ (.A(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__and2_1 _07058_ (.A(_06369_),
    .B(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__nand4_2 _07059_ (.A(net6),
    .B(net7),
    .C(net254),
    .D(net255),
    .Y(_06373_));
 sky130_fd_sc_hd__a21o_1 _07060_ (.A1(_05914_),
    .A2(_03787_),
    .B1(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_4 _07061_ (.A(net255),
    .X(_06375_));
 sky130_fd_sc_hd__a32o_1 _07062_ (.A1(_03798_),
    .A2(_05914_),
    .A3(_03831_),
    .B1(_06375_),
    .B2(_02470_),
    .X(_06376_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(_06374_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__xor2_1 _07064_ (.A(_06372_),
    .B(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__o21bai_1 _07065_ (.A1(_05893_),
    .A2(_05947_),
    .B1_N(_05936_),
    .Y(_06379_));
 sky130_fd_sc_hd__and2b_1 _07066_ (.A_N(_06378_),
    .B(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__and2b_1 _07067_ (.A_N(_06379_),
    .B(_06378_),
    .X(_06381_));
 sky130_fd_sc_hd__nor2_1 _07068_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__clkbuf_4 _07069_ (.A(net247),
    .X(_06383_));
 sky130_fd_sc_hd__buf_4 _07070_ (.A(net238),
    .X(_06384_));
 sky130_fd_sc_hd__and3_1 _07071_ (.A(net243),
    .B(net244),
    .C(net237),
    .X(_06385_));
 sky130_fd_sc_hd__a22o_1 _07072_ (.A1(net244),
    .A2(net237),
    .B1(net238),
    .B2(net243),
    .X(_06386_));
 sky130_fd_sc_hd__a21bo_1 _07073_ (.A1(_06384_),
    .A2(_06385_),
    .B1_N(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__nand2_1 _07074_ (.A(_03853_),
    .B(_05969_),
    .Y(_06388_));
 sky130_fd_sc_hd__xnor2_1 _07075_ (.A(_06387_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__a32o_1 _07076_ (.A1(net235),
    .A2(_05969_),
    .A3(_06001_),
    .B1(_03886_),
    .B2(_05980_),
    .X(_06390_));
 sky130_fd_sc_hd__xnor2_1 _07077_ (.A(_06389_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__and3_1 _07078_ (.A(_02503_),
    .B(_06383_),
    .C(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__a21oi_1 _07079_ (.A1(_02503_),
    .A2(_06383_),
    .B1(_06391_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _07080_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__xnor2_1 _07081_ (.A(_06382_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__nor2_1 _07082_ (.A(_06367_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__and2_1 _07083_ (.A(_06367_),
    .B(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__nor2_1 _07084_ (.A(_06396_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__and2_1 _07085_ (.A(_06366_),
    .B(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__nor2_1 _07086_ (.A(_06366_),
    .B(_06398_),
    .Y(_06400_));
 sky130_fd_sc_hd__or2_2 _07087_ (.A(_06399_),
    .B(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__or3_4 _07088_ (.A(_06359_),
    .B(_06360_),
    .C(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__o21ai_2 _07089_ (.A1(_06359_),
    .A2(_06360_),
    .B1(_06401_),
    .Y(_06403_));
 sky130_fd_sc_hd__o211ai_4 _07090_ (.A1(_05619_),
    .A2(_05663_),
    .B1(_06402_),
    .C1(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__a211o_1 _07091_ (.A1(_06402_),
    .A2(_06403_),
    .B1(_05619_),
    .C1(_05663_),
    .X(_06405_));
 sky130_fd_sc_hd__nand3_2 _07092_ (.A(_06112_),
    .B(_06404_),
    .C(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__a21o_1 _07093_ (.A1(_06404_),
    .A2(_06405_),
    .B1(_06112_),
    .X(_06407_));
 sky130_fd_sc_hd__inv_2 _07094_ (.A(_05356_),
    .Y(_06408_));
 sky130_fd_sc_hd__inv_2 _07095_ (.A(_05290_),
    .Y(_06409_));
 sky130_fd_sc_hd__buf_2 _07096_ (.A(net80),
    .X(_06410_));
 sky130_fd_sc_hd__or2_1 _07097_ (.A(_05487_),
    .B(_05531_),
    .X(_06411_));
 sky130_fd_sc_hd__and3_1 _07098_ (.A(_02668_),
    .B(_06410_),
    .C(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__a21oi_1 _07099_ (.A1(_02668_),
    .A2(_06410_),
    .B1(_06411_),
    .Y(_06413_));
 sky130_fd_sc_hd__nor2_1 _07100_ (.A(_06412_),
    .B(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__or3_1 _07101_ (.A(_05477_),
    .B(_05531_),
    .C(_05553_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_4 _07102_ (.A(net116),
    .X(_06416_));
 sky130_fd_sc_hd__a22o_1 _07103_ (.A1(net104),
    .A2(_05444_),
    .B1(_06416_),
    .B2(net103),
    .X(_06417_));
 sky130_fd_sc_hd__nand4_1 _07104_ (.A(net104),
    .B(net103),
    .C(_05444_),
    .D(_06416_),
    .Y(_06418_));
 sky130_fd_sc_hd__and3_1 _07105_ (.A(_05411_),
    .B(_06417_),
    .C(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__a21oi_1 _07106_ (.A1(_06417_),
    .A2(_06418_),
    .B1(_05411_),
    .Y(_06420_));
 sky130_fd_sc_hd__nor3_1 _07107_ (.A(_05455_),
    .B(_06419_),
    .C(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__o21a_1 _07108_ (.A1(_06419_),
    .A2(_06420_),
    .B1(_05455_),
    .X(_06422_));
 sky130_fd_sc_hd__and4_1 _07109_ (.A(net76),
    .B(net77),
    .C(net70),
    .D(net71),
    .X(_06423_));
 sky130_fd_sc_hd__clkbuf_4 _07110_ (.A(net71),
    .X(_06424_));
 sky130_fd_sc_hd__a22o_1 _07111_ (.A1(net77),
    .A2(_05498_),
    .B1(_06424_),
    .B2(net76),
    .X(_06425_));
 sky130_fd_sc_hd__or2b_1 _07112_ (.A(_06423_),
    .B_N(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__nand2_1 _07113_ (.A(_03579_),
    .B(_05520_),
    .Y(_06427_));
 sky130_fd_sc_hd__xnor2_1 _07114_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__or3_1 _07115_ (.A(_06421_),
    .B(_06422_),
    .C(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__o21ai_1 _07116_ (.A1(_06421_),
    .A2(_06422_),
    .B1(_06428_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(_06429_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__xor2_1 _07118_ (.A(_06415_),
    .B(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__nand2_1 _07119_ (.A(_06414_),
    .B(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__inv_2 _07120_ (.A(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__nor2_1 _07121_ (.A(_06414_),
    .B(_06432_),
    .Y(_06435_));
 sky130_fd_sc_hd__nor2_1 _07122_ (.A(_03425_),
    .B(_05422_),
    .Y(_06436_));
 sky130_fd_sc_hd__clkbuf_4 _07123_ (.A(net106),
    .X(_06437_));
 sky130_fd_sc_hd__a22o_1 _07124_ (.A1(_03546_),
    .A2(_05389_),
    .B1(_06437_),
    .B2(_02635_),
    .X(_00028_));
 sky130_fd_sc_hd__inv_2 _07125_ (.A(_00028_),
    .Y(_00029_));
 sky130_fd_sc_hd__and4_2 _07126_ (.A(_02635_),
    .B(_03546_),
    .C(_05389_),
    .D(_06437_),
    .X(_00030_));
 sky130_fd_sc_hd__or3_1 _07127_ (.A(_05246_),
    .B(_00029_),
    .C(_00030_),
    .X(_00031_));
 sky130_fd_sc_hd__o21ai_1 _07128_ (.A1(_00029_),
    .A2(_00030_),
    .B1(_05246_),
    .Y(_00032_));
 sky130_fd_sc_hd__and2_1 _07129_ (.A(_00031_),
    .B(_00032_),
    .X(_00033_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(_06436_),
    .B(_00033_),
    .Y(_00034_));
 sky130_fd_sc_hd__or2_1 _07131_ (.A(_06436_),
    .B(_00033_),
    .X(_00035_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(_00034_),
    .B(_00035_),
    .Y(_00036_));
 sky130_fd_sc_hd__or3_1 _07133_ (.A(_06434_),
    .B(_06435_),
    .C(_00036_),
    .X(_00037_));
 sky130_fd_sc_hd__o21ai_1 _07134_ (.A1(_06434_),
    .A2(_06435_),
    .B1(_00036_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _07135_ (.A(_00037_),
    .B(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__xnor2_1 _07136_ (.A(_06409_),
    .B(_00039_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _07137_ (.A(_05597_),
    .B(_00040_),
    .Y(_00041_));
 sky130_fd_sc_hd__or2_1 _07138_ (.A(_05597_),
    .B(_00040_),
    .X(_00042_));
 sky130_fd_sc_hd__and2_1 _07139_ (.A(_00041_),
    .B(_00042_),
    .X(_00043_));
 sky130_fd_sc_hd__or2b_1 _07140_ (.A(_04730_),
    .B_N(_05060_),
    .X(_00044_));
 sky130_fd_sc_hd__nor2_1 _07141_ (.A(_05180_),
    .B(_05268_),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _07142_ (.A(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__buf_2 _07143_ (.A(net185),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _07144_ (.A1(_03348_),
    .A2(net184),
    .B1(_00047_),
    .B2(net191),
    .X(_00048_));
 sky130_fd_sc_hd__buf_2 _07145_ (.A(_00047_),
    .X(_00049_));
 sky130_fd_sc_hd__nand4_1 _07146_ (.A(_02712_),
    .B(_03348_),
    .C(_05115_),
    .D(_00049_),
    .Y(_00050_));
 sky130_fd_sc_hd__a22oi_2 _07147_ (.A1(_03337_),
    .A2(_05093_),
    .B1(_00048_),
    .B2(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__and4_1 _07148_ (.A(_03337_),
    .B(_05093_),
    .C(_00048_),
    .D(_00050_),
    .X(_00052_));
 sky130_fd_sc_hd__a211o_1 _07149_ (.A1(_05126_),
    .A2(_05147_),
    .B1(_00051_),
    .C1(_00052_),
    .X(_00053_));
 sky130_fd_sc_hd__o211ai_1 _07150_ (.A1(_00051_),
    .A2(_00052_),
    .B1(_05126_),
    .C1(_05147_),
    .Y(_00054_));
 sky130_fd_sc_hd__and3_1 _07151_ (.A(_05158_),
    .B(_00053_),
    .C(_00054_),
    .X(_00055_));
 sky130_fd_sc_hd__a21oi_1 _07152_ (.A1(_00053_),
    .A2(_00054_),
    .B1(_05158_),
    .Y(_00056_));
 sky130_fd_sc_hd__nor2_1 _07153_ (.A(_00055_),
    .B(_00056_),
    .Y(_00057_));
 sky130_fd_sc_hd__clkbuf_4 _07154_ (.A(net194),
    .X(_00058_));
 sky130_fd_sc_hd__clkbuf_4 _07155_ (.A(net111),
    .X(_00059_));
 sky130_fd_sc_hd__a22oi_2 _07156_ (.A1(_02723_),
    .A2(_00058_),
    .B1(_00059_),
    .B2(_02734_),
    .Y(_00060_));
 sky130_fd_sc_hd__and4_1 _07157_ (.A(_02723_),
    .B(_02734_),
    .C(_00058_),
    .D(_00059_),
    .X(_00061_));
 sky130_fd_sc_hd__buf_2 _07158_ (.A(net176),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _07159_ (.A1(_03392_),
    .A2(_05191_),
    .B1(_05202_),
    .B2(_03381_),
    .X(_00063_));
 sky130_fd_sc_hd__nand4_4 _07160_ (.A(_03381_),
    .B(_03392_),
    .C(_05191_),
    .D(_05202_),
    .Y(_00064_));
 sky130_fd_sc_hd__a22o_1 _07161_ (.A1(_02745_),
    .A2(_00062_),
    .B1(_00063_),
    .B2(_00064_),
    .X(_00065_));
 sky130_fd_sc_hd__nand4_2 _07162_ (.A(_02745_),
    .B(_00062_),
    .C(_00063_),
    .D(_00064_),
    .Y(_00066_));
 sky130_fd_sc_hd__and3_1 _07163_ (.A(_05224_),
    .B(_00065_),
    .C(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__a21oi_1 _07164_ (.A1(_00065_),
    .A2(_00066_),
    .B1(_05224_),
    .Y(_00068_));
 sky130_fd_sc_hd__nor4_1 _07165_ (.A(_00060_),
    .B(_00061_),
    .C(_00067_),
    .D(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__o22a_1 _07166_ (.A1(_00060_),
    .A2(_00061_),
    .B1(_00067_),
    .B2(_00068_),
    .X(_00070_));
 sky130_fd_sc_hd__nor2_1 _07167_ (.A(_00069_),
    .B(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(_00057_),
    .B(_00071_),
    .Y(_00072_));
 sky130_fd_sc_hd__or2_1 _07169_ (.A(_00057_),
    .B(_00071_),
    .X(_00073_));
 sky130_fd_sc_hd__nand2_1 _07170_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__nor2_1 _07171_ (.A(_00046_),
    .B(_00074_),
    .Y(_00075_));
 sky130_fd_sc_hd__and2_1 _07172_ (.A(_00046_),
    .B(_00074_),
    .X(_00076_));
 sky130_fd_sc_hd__or2_1 _07173_ (.A(_00075_),
    .B(_00076_),
    .X(_00077_));
 sky130_fd_sc_hd__and2b_1 _07174_ (.A_N(_05016_),
    .B(_05038_),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _07175_ (.A(_04851_),
    .B(_05049_),
    .X(_00079_));
 sky130_fd_sc_hd__clkbuf_4 _07176_ (.A(net220),
    .X(_00080_));
 sky130_fd_sc_hd__and4_1 _07177_ (.A(net226),
    .B(_03260_),
    .C(_04752_),
    .D(_00080_),
    .X(_00081_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(_03227_),
    .B(_02855_),
    .Y(_00082_));
 sky130_fd_sc_hd__a32o_1 _07179_ (.A1(_03260_),
    .A2(_04752_),
    .A3(_00082_),
    .B1(_00080_),
    .B2(_02855_),
    .X(_00083_));
 sky130_fd_sc_hd__a21bo_1 _07180_ (.A1(_04785_),
    .A2(_00081_),
    .B1_N(_00083_),
    .X(_00084_));
 sky130_fd_sc_hd__xor2_1 _07181_ (.A(_04796_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__clkbuf_4 _07182_ (.A(net229),
    .X(_00086_));
 sky130_fd_sc_hd__a22oi_1 _07183_ (.A1(_03227_),
    .A2(_04741_),
    .B1(_00086_),
    .B2(_02866_),
    .Y(_00087_));
 sky130_fd_sc_hd__and4_1 _07184_ (.A(_03227_),
    .B(_02866_),
    .C(_04741_),
    .D(_00086_),
    .X(_00088_));
 sky130_fd_sc_hd__nor2_1 _07185_ (.A(_00087_),
    .B(_00088_),
    .Y(_00089_));
 sky130_fd_sc_hd__and2_1 _07186_ (.A(_00085_),
    .B(_00089_),
    .X(_00090_));
 sky130_fd_sc_hd__nor2_1 _07187_ (.A(_00085_),
    .B(_00089_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor2_1 _07188_ (.A(_00090_),
    .B(_00091_),
    .Y(_00092_));
 sky130_fd_sc_hd__and2_1 _07189_ (.A(_04818_),
    .B(_00092_),
    .X(_00093_));
 sky130_fd_sc_hd__nor2_1 _07190_ (.A(_04818_),
    .B(_00092_),
    .Y(_00094_));
 sky130_fd_sc_hd__or2_1 _07191_ (.A(_00093_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__and4_1 _07192_ (.A(net33),
    .B(net42),
    .C(net35),
    .D(net43),
    .X(_00096_));
 sky130_fd_sc_hd__buf_2 _07193_ (.A(net44),
    .X(_00097_));
 sky130_fd_sc_hd__a22o_1 _07194_ (.A1(net42),
    .A2(net35),
    .B1(net43),
    .B2(net33),
    .X(_00098_));
 sky130_fd_sc_hd__and4b_1 _07195_ (.A_N(_00096_),
    .B(_00097_),
    .C(net32),
    .D(_00098_),
    .X(_00099_));
 sky130_fd_sc_hd__inv_2 _07196_ (.A(_00096_),
    .Y(_00100_));
 sky130_fd_sc_hd__a22oi_1 _07197_ (.A1(_02822_),
    .A2(_00097_),
    .B1(_00098_),
    .B2(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__nor2_1 _07198_ (.A(_00099_),
    .B(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__and2_1 _07199_ (.A(_04884_),
    .B(_00102_),
    .X(_00103_));
 sky130_fd_sc_hd__nor2_1 _07200_ (.A(_04884_),
    .B(_00102_),
    .Y(_00104_));
 sky130_fd_sc_hd__or2_1 _07201_ (.A(_00103_),
    .B(_00104_),
    .X(_00105_));
 sky130_fd_sc_hd__and3_1 _07202_ (.A(_02811_),
    .B(_04906_),
    .C(_04983_),
    .X(_00106_));
 sky130_fd_sc_hd__clkbuf_4 _07203_ (.A(net36),
    .X(_00107_));
 sky130_fd_sc_hd__and3_1 _07204_ (.A(_02800_),
    .B(_03128_),
    .C(_04972_),
    .X(_00108_));
 sky130_fd_sc_hd__buf_2 _07205_ (.A(net23),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _07206_ (.A(_02800_),
    .B(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__and2_1 _07207_ (.A(net112),
    .B(net12),
    .X(_00111_));
 sky130_fd_sc_hd__nand4_1 _07208_ (.A(net245),
    .B(net256),
    .C(net179),
    .D(net190),
    .Y(_00112_));
 sky130_fd_sc_hd__a22o_1 _07209_ (.A1(net256),
    .A2(net179),
    .B1(net190),
    .B2(net245),
    .X(_00113_));
 sky130_fd_sc_hd__nand3_1 _07210_ (.A(_00111_),
    .B(_00112_),
    .C(_00113_),
    .Y(_00114_));
 sky130_fd_sc_hd__a21o_1 _07211_ (.A1(_00112_),
    .A2(_00113_),
    .B1(_00111_),
    .X(_00115_));
 sky130_fd_sc_hd__a32o_1 _07212_ (.A1(net1),
    .A2(net12),
    .A3(_04950_),
    .B1(_03128_),
    .B2(_04939_),
    .X(_00116_));
 sky130_fd_sc_hd__and3_1 _07213_ (.A(_00114_),
    .B(_00115_),
    .C(_00116_),
    .X(_00117_));
 sky130_fd_sc_hd__a21oi_2 _07214_ (.A1(_00114_),
    .A2(_00115_),
    .B1(net316),
    .Y(_00118_));
 sky130_fd_sc_hd__or3_4 _07215_ (.A(_00110_),
    .B(_00117_),
    .C(_00118_),
    .X(_00119_));
 sky130_fd_sc_hd__o21ai_1 _07216_ (.A1(net315),
    .A2(_00118_),
    .B1(_00110_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand3_1 _07217_ (.A(_00108_),
    .B(net317),
    .C(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__a21o_1 _07218_ (.A1(_00119_),
    .A2(_00120_),
    .B1(_00108_),
    .X(_00122_));
 sky130_fd_sc_hd__nand4_2 _07219_ (.A(_02811_),
    .B(_00107_),
    .C(_00121_),
    .D(_00122_),
    .Y(_00123_));
 sky130_fd_sc_hd__a22o_1 _07220_ (.A1(_02811_),
    .A2(_00107_),
    .B1(_00121_),
    .B2(_00122_),
    .X(_00124_));
 sky130_fd_sc_hd__and3_1 _07221_ (.A(_00106_),
    .B(_00123_),
    .C(_00124_),
    .X(_00125_));
 sky130_fd_sc_hd__a21oi_1 _07222_ (.A1(_00123_),
    .A2(_00124_),
    .B1(_00106_),
    .Y(_00126_));
 sky130_fd_sc_hd__or3_4 _07223_ (.A(_00105_),
    .B(_00125_),
    .C(_00126_),
    .X(_00127_));
 sky130_fd_sc_hd__o21ai_1 _07224_ (.A1(_00125_),
    .A2(_00126_),
    .B1(_00105_),
    .Y(_00128_));
 sky130_fd_sc_hd__and2_1 _07225_ (.A(_03150_),
    .B(_04994_),
    .X(_00129_));
 sky130_fd_sc_hd__a21o_1 _07226_ (.A1(_04895_),
    .A2(_05005_),
    .B1(_00129_),
    .X(_00130_));
 sky130_fd_sc_hd__and3_4 _07227_ (.A(_00127_),
    .B(_00128_),
    .C(_00130_),
    .X(_00131_));
 sky130_fd_sc_hd__a21oi_2 _07228_ (.A1(_00127_),
    .A2(_00128_),
    .B1(_00130_),
    .Y(_00132_));
 sky130_fd_sc_hd__or3_4 _07229_ (.A(_00095_),
    .B(_00131_),
    .C(_00132_),
    .X(_00133_));
 sky130_fd_sc_hd__o21ai_1 _07230_ (.A1(_00131_),
    .A2(_00132_),
    .B1(_00095_),
    .Y(_00134_));
 sky130_fd_sc_hd__o211a_2 _07231_ (.A1(_00078_),
    .A2(_00079_),
    .B1(_00133_),
    .C1(_00134_),
    .X(_00135_));
 sky130_fd_sc_hd__a211oi_4 _07232_ (.A1(_00133_),
    .A2(_00134_),
    .B1(_00078_),
    .C1(_00079_),
    .Y(_00136_));
 sky130_fd_sc_hd__nor3_2 _07233_ (.A(_00077_),
    .B(_00135_),
    .C(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__o21a_1 _07234_ (.A1(_00135_),
    .A2(_00136_),
    .B1(_00077_),
    .X(_00138_));
 sky130_fd_sc_hd__a211o_1 _07235_ (.A1(_00044_),
    .A2(_05323_),
    .B1(_00137_),
    .C1(_00138_),
    .X(_00139_));
 sky130_fd_sc_hd__o211ai_2 _07236_ (.A1(_00137_),
    .A2(_00138_),
    .B1(_00044_),
    .C1(_05323_),
    .Y(_00140_));
 sky130_fd_sc_hd__and3_2 _07237_ (.A(_00043_),
    .B(_00139_),
    .C(_00140_),
    .X(_00141_));
 sky130_fd_sc_hd__a21oi_1 _07238_ (.A1(_00139_),
    .A2(_00140_),
    .B1(_00043_),
    .Y(_00142_));
 sky130_fd_sc_hd__a211o_1 _07239_ (.A1(_06408_),
    .A2(_05696_),
    .B1(_00141_),
    .C1(_00142_),
    .X(_00143_));
 sky130_fd_sc_hd__o211ai_2 _07240_ (.A1(_00141_),
    .A2(_00142_),
    .B1(_06408_),
    .C1(_05696_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand4_2 _07241_ (.A(_06406_),
    .B(_06407_),
    .C(_00143_),
    .D(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__a22o_1 _07242_ (.A1(_06406_),
    .A2(_06407_),
    .B1(_00143_),
    .B2(_00144_),
    .X(_00146_));
 sky130_fd_sc_hd__o211a_2 _07243_ (.A1(_05729_),
    .A2(_06341_),
    .B1(_00145_),
    .C1(_00146_),
    .X(_00147_));
 sky130_fd_sc_hd__a211oi_1 _07244_ (.A1(_00145_),
    .A2(_00146_),
    .B1(_05729_),
    .C1(_06341_),
    .Y(_00148_));
 sky130_fd_sc_hd__nor4_1 _07245_ (.A(_06339_),
    .B(_06340_),
    .C(_00147_),
    .D(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__o22a_1 _07246_ (.A1(_06339_),
    .A2(_06340_),
    .B1(_00147_),
    .B2(_00148_),
    .X(_00150_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(_06125_),
    .B(_06203_),
    .Y(_00151_));
 sky130_fd_sc_hd__or3_2 _07248_ (.A(_00149_),
    .B(_00150_),
    .C(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__o21ai_1 _07249_ (.A1(_00149_),
    .A2(_00150_),
    .B1(_00151_),
    .Y(_00153_));
 sky130_fd_sc_hd__and3_2 _07250_ (.A(_06241_),
    .B(_00152_),
    .C(_00153_),
    .X(_00154_));
 sky130_fd_sc_hd__a21oi_2 _07251_ (.A1(_00152_),
    .A2(_00153_),
    .B1(_06241_),
    .Y(_00155_));
 sky130_fd_sc_hd__a211oi_4 _07252_ (.A1(_06225_),
    .A2(_06214_),
    .B1(_00154_),
    .C1(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__o211a_1 _07253_ (.A1(_00154_),
    .A2(_00155_),
    .B1(_06225_),
    .C1(_06214_),
    .X(_00157_));
 sky130_fd_sc_hd__or3_1 _07254_ (.A(_06211_),
    .B(_00156_),
    .C(_00157_),
    .X(_00158_));
 sky130_fd_sc_hd__o21ai_2 _07255_ (.A1(_00156_),
    .A2(_00157_),
    .B1(_06211_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand3_2 _07256_ (.A(_06224_),
    .B(_00158_),
    .C(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__a21o_1 _07257_ (.A1(_00158_),
    .A2(_00159_),
    .B1(_06224_),
    .X(_00161_));
 sky130_fd_sc_hd__nand3_1 _07258_ (.A(net279),
    .B(_00160_),
    .C(_00161_),
    .Y(_00162_));
 sky130_fd_sc_hd__a21o_1 _07259_ (.A1(_00160_),
    .A2(_00161_),
    .B1(net279),
    .X(_00163_));
 sky130_fd_sc_hd__a21bo_1 _07260_ (.A1(net278),
    .A2(_06218_),
    .B1_N(_06222_),
    .X(_00164_));
 sky130_fd_sc_hd__a21oi_1 _07261_ (.A1(_00162_),
    .A2(_00163_),
    .B1(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__clkinv_4 _07262_ (.A(net257),
    .Y(_00166_));
 sky130_fd_sc_hd__a31o_1 _07263_ (.A1(_00162_),
    .A2(_00163_),
    .A3(_00164_),
    .B1(_00166_),
    .X(_00167_));
 sky130_fd_sc_hd__nor2_1 _07264_ (.A(_00165_),
    .B(_00167_),
    .Y(_00003_));
 sky130_fd_sc_hd__nor3_1 _07265_ (.A(_06211_),
    .B(_00156_),
    .C(_00157_),
    .Y(_00168_));
 sky130_fd_sc_hd__inv_2 _07266_ (.A(_00152_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_06226_),
    .B(_06234_),
    .Y(_00170_));
 sky130_fd_sc_hd__clkbuf_4 _07268_ (.A(net170),
    .X(_00171_));
 sky130_fd_sc_hd__nand4_1 _07269_ (.A(_04227_),
    .B(_02328_),
    .C(_06227_),
    .D(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__a22o_1 _07270_ (.A1(_04227_),
    .A2(_06227_),
    .B1(_00171_),
    .B2(net157),
    .X(_00173_));
 sky130_fd_sc_hd__and2_1 _07271_ (.A(_00172_),
    .B(_00173_),
    .X(_00174_));
 sky130_fd_sc_hd__o21ai_1 _07272_ (.A1(_06245_),
    .A2(_06248_),
    .B1(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__or3_1 _07273_ (.A(_06245_),
    .B(_06248_),
    .C(_00174_),
    .X(_00176_));
 sky130_fd_sc_hd__and2_1 _07274_ (.A(_00175_),
    .B(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__nand2_1 _07275_ (.A(_06229_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__or2_1 _07276_ (.A(_06229_),
    .B(_00177_),
    .X(_00179_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(_00178_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__nor3_1 _07278_ (.A(_06148_),
    .B(_06251_),
    .C(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__o21a_1 _07279_ (.A1(_06148_),
    .A2(_06251_),
    .B1(_00180_),
    .X(_00182_));
 sky130_fd_sc_hd__or2_1 _07280_ (.A(net303),
    .B(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__a21bo_1 _07281_ (.A1(_06252_),
    .A2(_06298_),
    .B1_N(_06297_),
    .X(_00184_));
 sky130_fd_sc_hd__and2b_1 _07282_ (.A_N(_00183_),
    .B(_00184_),
    .X(_00185_));
 sky130_fd_sc_hd__and2b_1 _07283_ (.A_N(_00184_),
    .B(_00183_),
    .X(_00186_));
 sky130_fd_sc_hd__nor2_1 _07284_ (.A(_00185_),
    .B(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__xor2_1 _07285_ (.A(_06232_),
    .B(_00187_),
    .X(_00188_));
 sky130_fd_sc_hd__o21a_1 _07286_ (.A1(_06337_),
    .A2(_06339_),
    .B1(_00188_),
    .X(_00189_));
 sky130_fd_sc_hd__nor3_1 _07287_ (.A(_06337_),
    .B(_06339_),
    .C(_00188_),
    .Y(_00190_));
 sky130_fd_sc_hd__nor2_1 _07288_ (.A(_00189_),
    .B(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__xnor2_1 _07289_ (.A(_00170_),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__or2_1 _07290_ (.A(_06189_),
    .B(_06333_),
    .X(_00193_));
 sky130_fd_sc_hd__nand2_1 _07291_ (.A(_06301_),
    .B(_06335_),
    .Y(_00194_));
 sky130_fd_sc_hd__or3b_1 _07292_ (.A(_04358_),
    .B(_06161_),
    .C_N(_06288_),
    .X(_00195_));
 sky130_fd_sc_hd__or2b_1 _07293_ (.A(_06289_),
    .B_N(_06288_),
    .X(_00196_));
 sky130_fd_sc_hd__inv_2 _07294_ (.A(_06273_),
    .Y(_00197_));
 sky130_fd_sc_hd__nor2_1 _07295_ (.A(_00197_),
    .B(_06281_),
    .Y(_00198_));
 sky130_fd_sc_hd__and2b_1 _07296_ (.A_N(_06282_),
    .B(_06287_),
    .X(_00199_));
 sky130_fd_sc_hd__clkbuf_4 _07297_ (.A(net90),
    .X(_00200_));
 sky130_fd_sc_hd__buf_2 _07298_ (.A(net135),
    .X(_00201_));
 sky130_fd_sc_hd__a22o_1 _07299_ (.A1(_04303_),
    .A2(_06283_),
    .B1(_00201_),
    .B2(_02229_),
    .X(_00202_));
 sky130_fd_sc_hd__and4_1 _07300_ (.A(net122),
    .B(net121),
    .C(_06283_),
    .D(_00201_),
    .X(_00203_));
 sky130_fd_sc_hd__inv_2 _07301_ (.A(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand4_2 _07302_ (.A(_02240_),
    .B(_00200_),
    .C(_00202_),
    .D(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__a22o_1 _07303_ (.A1(_02240_),
    .A2(_00200_),
    .B1(_00202_),
    .B2(_00204_),
    .X(_00206_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(_00205_),
    .B(_00206_),
    .Y(_00207_));
 sky130_fd_sc_hd__or2b_1 _07305_ (.A(_06279_),
    .B_N(_06280_),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_1 _07306_ (.A1(net131),
    .A2(net125),
    .B1(net126),
    .B2(net130),
    .X(_00209_));
 sky130_fd_sc_hd__buf_2 _07307_ (.A(net126),
    .X(_00210_));
 sky130_fd_sc_hd__nand4_1 _07308_ (.A(net130),
    .B(net131),
    .C(net125),
    .D(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__a22oi_1 _07309_ (.A1(_06152_),
    .A2(_06151_),
    .B1(_00209_),
    .B2(_00211_),
    .Y(_00212_));
 sky130_fd_sc_hd__and4_1 _07310_ (.A(net124),
    .B(net132),
    .C(_00209_),
    .D(_00211_),
    .X(_00213_));
 sky130_fd_sc_hd__a21bo_1 _07311_ (.A1(_06276_),
    .A2(_06278_),
    .B1_N(_06275_),
    .X(_00214_));
 sky130_fd_sc_hd__or3b_2 _07312_ (.A(_00212_),
    .B(_00213_),
    .C_N(_00214_),
    .X(_00215_));
 sky130_fd_sc_hd__o21bai_1 _07313_ (.A1(_00212_),
    .A2(_00213_),
    .B1_N(_00214_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _07314_ (.A(_00215_),
    .B(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__xnor2_1 _07315_ (.A(_00208_),
    .B(_00217_),
    .Y(_00218_));
 sky130_fd_sc_hd__xor2_1 _07316_ (.A(_00207_),
    .B(_00218_),
    .X(_00219_));
 sky130_fd_sc_hd__xor2_1 _07317_ (.A(_06323_),
    .B(_00219_),
    .X(_00220_));
 sky130_fd_sc_hd__o21a_1 _07318_ (.A1(_00198_),
    .A2(_00199_),
    .B1(_00220_),
    .X(_00221_));
 sky130_fd_sc_hd__nor3_1 _07319_ (.A(_00198_),
    .B(_00199_),
    .C(_00220_),
    .Y(_00222_));
 sky130_fd_sc_hd__or2_2 _07320_ (.A(_00221_),
    .B(_00222_),
    .X(_00223_));
 sky130_fd_sc_hd__xor2_1 _07321_ (.A(_00196_),
    .B(_00223_),
    .X(_00224_));
 sky130_fd_sc_hd__and2_1 _07322_ (.A(_06136_),
    .B(_06259_),
    .X(_00225_));
 sky130_fd_sc_hd__inv_2 _07323_ (.A(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__a22o_1 _07324_ (.A1(net87),
    .A2(_06254_),
    .B1(net88),
    .B2(_04413_),
    .X(_00227_));
 sky130_fd_sc_hd__nand4_1 _07325_ (.A(_04424_),
    .B(net87),
    .C(_06134_),
    .D(net88),
    .Y(_00228_));
 sky130_fd_sc_hd__a22oi_1 _07326_ (.A1(_04292_),
    .A2(_06253_),
    .B1(_00227_),
    .B2(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__and4_1 _07327_ (.A(net86),
    .B(_06253_),
    .C(_00227_),
    .D(_00228_),
    .X(_00230_));
 sky130_fd_sc_hd__nor2_1 _07328_ (.A(_00229_),
    .B(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__a41o_1 _07329_ (.A1(_04292_),
    .A2(_04424_),
    .A3(_06159_),
    .A4(_06134_),
    .B1(_06257_),
    .X(_00232_));
 sky130_fd_sc_hd__xnor2_2 _07330_ (.A(_00231_),
    .B(_00232_),
    .Y(_00233_));
 sky130_fd_sc_hd__xnor2_1 _07331_ (.A(_06286_),
    .B(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__or2_1 _07332_ (.A(_00226_),
    .B(_00234_),
    .X(_00235_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(_00226_),
    .B(_00234_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _07334_ (.A(_00235_),
    .B(_00236_),
    .Y(_00237_));
 sky130_fd_sc_hd__clkbuf_4 _07335_ (.A(net98),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_4 _07336_ (.A(net19),
    .X(_00239_));
 sky130_fd_sc_hd__a22o_1 _07337_ (.A1(net25),
    .A2(_06261_),
    .B1(_00239_),
    .B2(net24),
    .X(_00240_));
 sky130_fd_sc_hd__nand4_2 _07338_ (.A(_02196_),
    .B(_04446_),
    .C(_06261_),
    .D(_00239_),
    .Y(_00241_));
 sky130_fd_sc_hd__and4_1 _07339_ (.A(_02251_),
    .B(_00238_),
    .C(_00240_),
    .D(_00241_),
    .X(_00242_));
 sky130_fd_sc_hd__inv_2 _07340_ (.A(_00242_),
    .Y(_00243_));
 sky130_fd_sc_hd__a22o_1 _07341_ (.A1(_02251_),
    .A2(_00238_),
    .B1(_00240_),
    .B2(_00241_),
    .X(_00244_));
 sky130_fd_sc_hd__and2_1 _07342_ (.A(_00243_),
    .B(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__inv_2 _07343_ (.A(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__a22o_1 _07344_ (.A1(net17),
    .A2(net26),
    .B1(net27),
    .B2(net16),
    .X(_00247_));
 sky130_fd_sc_hd__nand4_1 _07345_ (.A(net16),
    .B(_06138_),
    .C(_06142_),
    .D(_06264_),
    .Y(_00248_));
 sky130_fd_sc_hd__a22o_1 _07346_ (.A1(net15),
    .A2(net28),
    .B1(_00247_),
    .B2(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__buf_2 _07347_ (.A(net28),
    .X(_00250_));
 sky130_fd_sc_hd__nand4_1 _07348_ (.A(net15),
    .B(_00250_),
    .C(_00247_),
    .D(_00248_),
    .Y(_00251_));
 sky130_fd_sc_hd__and3_1 _07349_ (.A(_06263_),
    .B(_00249_),
    .C(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__a21oi_1 _07350_ (.A1(_00249_),
    .A2(_00251_),
    .B1(_06263_),
    .Y(_00253_));
 sky130_fd_sc_hd__or2_1 _07351_ (.A(_00252_),
    .B(_00253_),
    .X(_00254_));
 sky130_fd_sc_hd__xnor2_1 _07352_ (.A(_06265_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(_00246_),
    .B(_00255_),
    .Y(_00256_));
 sky130_fd_sc_hd__and2_1 _07354_ (.A(_00246_),
    .B(_00255_),
    .X(_00257_));
 sky130_fd_sc_hd__or2_1 _07355_ (.A(_00256_),
    .B(_00257_),
    .X(_00258_));
 sky130_fd_sc_hd__or2_1 _07356_ (.A(_00237_),
    .B(_00258_),
    .X(_00259_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_00237_),
    .B(_00258_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(_00259_),
    .B(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _07359_ (.A(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__xnor2_1 _07360_ (.A(_00224_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__a21oi_2 _07361_ (.A1(_06292_),
    .A2(_00195_),
    .B1(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__and3_1 _07362_ (.A(_06292_),
    .B(_00263_),
    .C(_00195_),
    .X(_00265_));
 sky130_fd_sc_hd__or3_1 _07363_ (.A(_06260_),
    .B(_06269_),
    .C(_06270_),
    .X(_00266_));
 sky130_fd_sc_hd__inv_2 _07364_ (.A(_06142_),
    .Y(_00267_));
 sky130_fd_sc_hd__or4_1 _07365_ (.A(_00267_),
    .B(_04479_),
    .C(_06247_),
    .D(_06248_),
    .X(_00268_));
 sky130_fd_sc_hd__inv_2 _07366_ (.A(net308),
    .Y(_00269_));
 sky130_fd_sc_hd__clkbuf_4 _07367_ (.A(net161),
    .X(_00270_));
 sky130_fd_sc_hd__a22o_1 _07368_ (.A1(_04238_),
    .A2(_06243_),
    .B1(_00270_),
    .B2(_02317_),
    .X(_00271_));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__and4_1 _07370_ (.A(_02317_),
    .B(_04238_),
    .C(_06243_),
    .D(_00270_),
    .X(_00273_));
 sky130_fd_sc_hd__o2bb2a_1 _07371_ (.A1_N(_06127_),
    .A2_N(_06130_),
    .B1(_00272_),
    .B2(_00273_),
    .X(_00274_));
 sky130_fd_sc_hd__and4b_1 _07372_ (.A_N(_00273_),
    .B(_06130_),
    .C(_06127_),
    .D(_00271_),
    .X(_00275_));
 sky130_fd_sc_hd__or2_1 _07373_ (.A(_00274_),
    .B(_00275_),
    .X(_00276_));
 sky130_fd_sc_hd__or3b_1 _07374_ (.A(_06267_),
    .B(net308),
    .C_N(_00276_),
    .X(_00277_));
 sky130_fd_sc_hd__or3b_2 _07375_ (.A(_00274_),
    .B(_00275_),
    .C_N(_06267_),
    .X(_00278_));
 sky130_fd_sc_hd__o211a_1 _07376_ (.A1(_00269_),
    .A2(_00276_),
    .B1(_00277_),
    .C1(_00278_),
    .X(_00279_));
 sky130_fd_sc_hd__xor2_1 _07377_ (.A(_00268_),
    .B(_00279_),
    .X(_00280_));
 sky130_fd_sc_hd__nor2_1 _07378_ (.A(_00266_),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__and2_1 _07379_ (.A(_00266_),
    .B(_00280_),
    .X(_00282_));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_00281_),
    .B(_00282_),
    .Y(_00283_));
 sky130_fd_sc_hd__and3_1 _07381_ (.A(_06145_),
    .B(_06249_),
    .C(_00283_),
    .X(_00284_));
 sky130_fd_sc_hd__a21oi_1 _07382_ (.A1(_06145_),
    .A2(_06249_),
    .B1(_00283_),
    .Y(_00285_));
 sky130_fd_sc_hd__nor2_1 _07383_ (.A(_00284_),
    .B(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__nor3b_2 _07384_ (.A(_00264_),
    .B(_00265_),
    .C_N(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__o21ba_1 _07385_ (.A1(_00264_),
    .A2(_00265_),
    .B1_N(_00286_),
    .X(_00288_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(_06182_),
    .B(_06317_),
    .Y(_00289_));
 sky130_fd_sc_hd__or2_1 _07387_ (.A(_06310_),
    .B(_06316_),
    .X(_00290_));
 sky130_fd_sc_hd__clkbuf_4 _07388_ (.A(net143),
    .X(_00291_));
 sky130_fd_sc_hd__nand4_2 _07389_ (.A(_02383_),
    .B(_04139_),
    .C(_06311_),
    .D(_00291_),
    .Y(_00292_));
 sky130_fd_sc_hd__and2b_1 _07390_ (.A_N(_00292_),
    .B(_06312_),
    .X(_00293_));
 sky130_fd_sc_hd__a22oi_1 _07391_ (.A1(_04139_),
    .A2(_06311_),
    .B1(_00291_),
    .B2(_02383_),
    .Y(_00294_));
 sky130_fd_sc_hd__and2b_1 _07392_ (.A_N(_06312_),
    .B(_00292_),
    .X(_00295_));
 sky130_fd_sc_hd__or3_2 _07393_ (.A(_00293_),
    .B(_00294_),
    .C(_00295_),
    .X(_00296_));
 sky130_fd_sc_hd__buf_2 _07394_ (.A(net213),
    .X(_00297_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(_02459_),
    .B(_00297_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand4_1 _07396_ (.A(net209),
    .B(_06077_),
    .C(_06172_),
    .D(_06361_),
    .Y(_00299_));
 sky130_fd_sc_hd__a22o_1 _07397_ (.A1(_06077_),
    .A2(net210),
    .B1(net203),
    .B2(net209),
    .X(_00300_));
 sky130_fd_sc_hd__nand4_1 _07398_ (.A(_03941_),
    .B(_06304_),
    .C(_00299_),
    .D(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__a22o_1 _07399_ (.A1(net200),
    .A2(net211),
    .B1(_00299_),
    .B2(_00300_),
    .X(_00302_));
 sky130_fd_sc_hd__a32o_1 _07400_ (.A1(net199),
    .A2(net211),
    .A3(_06307_),
    .B1(_06306_),
    .B2(_06077_),
    .X(_00303_));
 sky130_fd_sc_hd__and3_1 _07401_ (.A(_00301_),
    .B(_00302_),
    .C(_00303_),
    .X(_00304_));
 sky130_fd_sc_hd__a21oi_1 _07402_ (.A1(_00301_),
    .A2(_00302_),
    .B1(_00303_),
    .Y(_00305_));
 sky130_fd_sc_hd__or3_1 _07403_ (.A(_00298_),
    .B(_00304_),
    .C(_00305_),
    .X(_00306_));
 sky130_fd_sc_hd__o21ai_1 _07404_ (.A1(_00304_),
    .A2(_00305_),
    .B1(_00298_),
    .Y(_00307_));
 sky130_fd_sc_hd__and2_1 _07405_ (.A(_06175_),
    .B(_06309_),
    .X(_00308_));
 sky130_fd_sc_hd__a21o_1 _07406_ (.A1(_00306_),
    .A2(_00307_),
    .B1(_00308_),
    .X(_00309_));
 sky130_fd_sc_hd__nand3_1 _07407_ (.A(_00308_),
    .B(_00306_),
    .C(_00307_),
    .Y(_00310_));
 sky130_fd_sc_hd__and3b_1 _07408_ (.A_N(_00296_),
    .B(_00309_),
    .C(_00310_),
    .X(_00311_));
 sky130_fd_sc_hd__a21boi_1 _07409_ (.A1(_00310_),
    .A2(_00309_),
    .B1_N(_00296_),
    .Y(_00312_));
 sky130_fd_sc_hd__nor2_1 _07410_ (.A(_00311_),
    .B(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__xnor2_1 _07411_ (.A(_00290_),
    .B(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand4_1 _07412_ (.A(net140),
    .B(_06177_),
    .C(net150),
    .D(net151),
    .Y(_00315_));
 sky130_fd_sc_hd__a22o_1 _07413_ (.A1(net141),
    .A2(net150),
    .B1(net151),
    .B2(net140),
    .X(_00316_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(net139),
    .B(net152),
    .X(_00317_));
 sky130_fd_sc_hd__nand3_1 _07415_ (.A(_00315_),
    .B(_00316_),
    .C(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__a21o_1 _07416_ (.A1(_00315_),
    .A2(_00316_),
    .B1(_00317_),
    .X(_00319_));
 sky130_fd_sc_hd__and3_1 _07417_ (.A(_06322_),
    .B(_00318_),
    .C(_00319_),
    .X(_00320_));
 sky130_fd_sc_hd__a21oi_1 _07418_ (.A1(_00318_),
    .A2(_00319_),
    .B1(_06322_),
    .Y(_00321_));
 sky130_fd_sc_hd__or2_1 _07419_ (.A(_00320_),
    .B(_00321_),
    .X(_00322_));
 sky130_fd_sc_hd__or2_2 _07420_ (.A(_06315_),
    .B(_00322_),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_1 _07421_ (.A(_06315_),
    .B(_00322_),
    .Y(_00324_));
 sky130_fd_sc_hd__and2_1 _07422_ (.A(_00323_),
    .B(_00324_),
    .X(_00325_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(_00314_),
    .B(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__a21o_2 _07424_ (.A1(_00289_),
    .A2(_06326_),
    .B1(_00326_),
    .X(_00327_));
 sky130_fd_sc_hd__nand3_2 _07425_ (.A(_00289_),
    .B(_06326_),
    .C(_00326_),
    .Y(_00328_));
 sky130_fd_sc_hd__a211oi_2 _07426_ (.A1(_00327_),
    .A2(_00328_),
    .B1(_06396_),
    .C1(_06399_),
    .Y(_00329_));
 sky130_fd_sc_hd__o211a_1 _07427_ (.A1(_06396_),
    .A2(_06399_),
    .B1(_00327_),
    .C1(_00328_),
    .X(_00330_));
 sky130_fd_sc_hd__or2_2 _07428_ (.A(_00329_),
    .B(_00330_),
    .X(_00331_));
 sky130_fd_sc_hd__and2b_2 _07429_ (.A_N(_06329_),
    .B(_06328_),
    .X(_00332_));
 sky130_fd_sc_hd__and2b_1 _07430_ (.A_N(_00332_),
    .B(_06331_),
    .X(_00333_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(_00331_),
    .B(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__nor3_1 _07432_ (.A(_00287_),
    .B(_00288_),
    .C(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__o21a_1 _07433_ (.A1(_00287_),
    .A2(_00288_),
    .B1(_00334_),
    .X(_00336_));
 sky130_fd_sc_hd__a211oi_2 _07434_ (.A1(_06404_),
    .A2(_06406_),
    .B1(_00335_),
    .C1(_00336_),
    .Y(_00337_));
 sky130_fd_sc_hd__o211a_1 _07435_ (.A1(_00335_),
    .A2(_00336_),
    .B1(_06404_),
    .C1(_06406_),
    .X(_00338_));
 sky130_fd_sc_hd__a211oi_2 _07436_ (.A1(_00193_),
    .A2(_00194_),
    .B1(_00337_),
    .C1(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__o211a_1 _07437_ (.A1(_00337_),
    .A2(_00338_),
    .B1(_00193_),
    .C1(_00194_),
    .X(_00340_));
 sky130_fd_sc_hd__or2_1 _07438_ (.A(_06409_),
    .B(_00039_),
    .X(_00341_));
 sky130_fd_sc_hd__and2b_1 _07439_ (.A_N(_06389_),
    .B(_06390_),
    .X(_00342_));
 sky130_fd_sc_hd__clkbuf_4 _07440_ (.A(net204),
    .X(_00343_));
 sky130_fd_sc_hd__nand2_1 _07441_ (.A(_02448_),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__o21ba_1 _07442_ (.A1(_00342_),
    .A2(_06392_),
    .B1_N(_00344_),
    .X(_00345_));
 sky130_fd_sc_hd__nor3b_1 _07443_ (.A(_00342_),
    .B(_06392_),
    .C_N(_00344_),
    .Y(_00346_));
 sky130_fd_sc_hd__or2_1 _07444_ (.A(_00345_),
    .B(_00346_),
    .X(_00347_));
 sky130_fd_sc_hd__xor2_1 _07445_ (.A(_06364_),
    .B(_00347_),
    .X(_00348_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(_06382_),
    .B(_06394_),
    .Y(_00349_));
 sky130_fd_sc_hd__and4_1 _07447_ (.A(net253),
    .B(net254),
    .C(net8),
    .D(net9),
    .X(_00350_));
 sky130_fd_sc_hd__a22o_1 _07448_ (.A1(net254),
    .A2(net8),
    .B1(net9),
    .B2(net253),
    .X(_00351_));
 sky130_fd_sc_hd__and2b_1 _07449_ (.A_N(_00350_),
    .B(_00351_),
    .X(_00352_));
 sky130_fd_sc_hd__nand2_1 _07450_ (.A(net252),
    .B(net10),
    .Y(_00353_));
 sky130_fd_sc_hd__xnor2_2 _07451_ (.A(_00352_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__and4_1 _07452_ (.A(net6),
    .B(net7),
    .C(net255),
    .D(net2),
    .X(_00355_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(_06373_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__buf_4 _07454_ (.A(net2),
    .X(_00357_));
 sky130_fd_sc_hd__a22o_1 _07455_ (.A1(_03798_),
    .A2(net255),
    .B1(_00357_),
    .B2(_02470_),
    .X(_00358_));
 sky130_fd_sc_hd__or2_1 _07456_ (.A(_06373_),
    .B(_00355_),
    .X(_00359_));
 sky130_fd_sc_hd__and3_1 _07457_ (.A(_00356_),
    .B(_00358_),
    .C(_00359_),
    .X(_00360_));
 sky130_fd_sc_hd__xor2_1 _07458_ (.A(_00354_),
    .B(_00360_),
    .X(_00361_));
 sky130_fd_sc_hd__and3_1 _07459_ (.A(_05914_),
    .B(_03787_),
    .C(_06373_),
    .X(_00362_));
 sky130_fd_sc_hd__a31oi_2 _07460_ (.A1(_06372_),
    .A2(_06374_),
    .A3(_06376_),
    .B1(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__xnor2_1 _07461_ (.A(_00361_),
    .B(_00363_),
    .Y(_00364_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(_06380_),
    .B(_00364_),
    .Y(_00365_));
 sky130_fd_sc_hd__clkbuf_4 _07463_ (.A(net248),
    .X(_00366_));
 sky130_fd_sc_hd__a22oi_1 _07464_ (.A1(_03853_),
    .A2(_06383_),
    .B1(_00366_),
    .B2(_02503_),
    .Y(_00367_));
 sky130_fd_sc_hd__and4_1 _07465_ (.A(_03853_),
    .B(net235),
    .C(_06383_),
    .D(_00366_),
    .X(_00368_));
 sky130_fd_sc_hd__nor2_1 _07466_ (.A(_00367_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__a22o_1 _07467_ (.A1(net244),
    .A2(net238),
    .B1(net239),
    .B2(net243),
    .X(_00370_));
 sky130_fd_sc_hd__nand4_4 _07468_ (.A(net243),
    .B(net244),
    .C(net238),
    .D(net239),
    .Y(_00371_));
 sky130_fd_sc_hd__nand4_2 _07469_ (.A(_05980_),
    .B(_05969_),
    .C(_00370_),
    .D(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__a22o_1 _07470_ (.A1(_05980_),
    .A2(net246),
    .B1(_00370_),
    .B2(_00371_),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _07471_ (.A(_00372_),
    .B(_00373_),
    .Y(_00374_));
 sky130_fd_sc_hd__a32o_1 _07472_ (.A1(_03853_),
    .A2(_05969_),
    .A3(_06386_),
    .B1(_06385_),
    .B2(_06384_),
    .X(_00375_));
 sky130_fd_sc_hd__xnor2_1 _07473_ (.A(_00374_),
    .B(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__xnor2_1 _07474_ (.A(_00369_),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__xnor2_1 _07475_ (.A(_06371_),
    .B(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__nor2_1 _07476_ (.A(_00365_),
    .B(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__and2_1 _07477_ (.A(_00365_),
    .B(_00378_),
    .X(_00380_));
 sky130_fd_sc_hd__or3_2 _07478_ (.A(_00349_),
    .B(_00379_),
    .C(_00380_),
    .X(_00381_));
 sky130_fd_sc_hd__o21ai_1 _07479_ (.A1(_00379_),
    .A2(_00380_),
    .B1(_00349_),
    .Y(_00382_));
 sky130_fd_sc_hd__and3_2 _07480_ (.A(_00348_),
    .B(_00381_),
    .C(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__a21oi_2 _07481_ (.A1(_00381_),
    .A2(_00382_),
    .B1(_00348_),
    .Y(_00384_));
 sky130_fd_sc_hd__or2_1 _07482_ (.A(_06415_),
    .B(_06431_),
    .X(_00385_));
 sky130_fd_sc_hd__and4b_1 _07483_ (.A_N(_06348_),
    .B(_06350_),
    .C(_02569_),
    .D(_06343_),
    .X(_00386_));
 sky130_fd_sc_hd__clkbuf_4 _07484_ (.A(net54),
    .X(_00387_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(net52),
    .A2(_05761_),
    .B1(net53),
    .B2(_03743_),
    .X(_00388_));
 sky130_fd_sc_hd__nand4_1 _07486_ (.A(_03743_),
    .B(_05750_),
    .C(_05761_),
    .D(_06343_),
    .Y(_00389_));
 sky130_fd_sc_hd__and2_1 _07487_ (.A(net51),
    .B(net62),
    .X(_00390_));
 sky130_fd_sc_hd__a21o_1 _07488_ (.A1(_00388_),
    .A2(_00389_),
    .B1(_00390_),
    .X(_00391_));
 sky130_fd_sc_hd__nand3_1 _07489_ (.A(_00388_),
    .B(_00389_),
    .C(_00390_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand4_2 _07490_ (.A(_02569_),
    .B(_00387_),
    .C(_00391_),
    .D(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__a22o_1 _07491_ (.A1(net59),
    .A2(_00387_),
    .B1(_00391_),
    .B2(_00392_),
    .X(_00394_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(_00393_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__xnor2_1 _07493_ (.A(_00386_),
    .B(_00395_),
    .Y(_00396_));
 sky130_fd_sc_hd__clkbuf_4 _07494_ (.A(net63),
    .X(_00397_));
 sky130_fd_sc_hd__o211a_1 _07495_ (.A1(_06345_),
    .A2(_06348_),
    .B1(_02580_),
    .C1(_00397_),
    .X(_00398_));
 sky130_fd_sc_hd__a211oi_1 _07496_ (.A1(_02580_),
    .A2(_00397_),
    .B1(_06345_),
    .C1(_06348_),
    .Y(_00399_));
 sky130_fd_sc_hd__nor2_1 _07497_ (.A(_00398_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__xnor2_1 _07498_ (.A(_00396_),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__o21a_1 _07499_ (.A1(_05783_),
    .A2(_05805_),
    .B1(_06352_),
    .X(_00402_));
 sky130_fd_sc_hd__nor2b_1 _07500_ (.A(_00401_),
    .B_N(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__and2b_1 _07501_ (.A_N(_00402_),
    .B(_00401_),
    .X(_00404_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(_00403_),
    .B(_00404_),
    .X(_00405_));
 sky130_fd_sc_hd__and3_1 _07503_ (.A(_00385_),
    .B(_06433_),
    .C(_00405_),
    .X(_00406_));
 sky130_fd_sc_hd__a21o_1 _07504_ (.A1(_00385_),
    .A2(_06433_),
    .B1(_00405_),
    .X(_00407_));
 sky130_fd_sc_hd__or2b_1 _07505_ (.A(_00406_),
    .B_N(_00407_),
    .X(_00408_));
 sky130_fd_sc_hd__inv_2 _07506_ (.A(_06357_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2_1 _07507_ (.A(_00409_),
    .B(_06359_),
    .Y(_00410_));
 sky130_fd_sc_hd__xnor2_1 _07508_ (.A(_00408_),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__nor3_1 _07509_ (.A(_00383_),
    .B(_00384_),
    .C(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__o21a_1 _07510_ (.A1(_00383_),
    .A2(_00384_),
    .B1(_00411_),
    .X(_00413_));
 sky130_fd_sc_hd__a211oi_2 _07511_ (.A1(_00341_),
    .A2(_00042_),
    .B1(net296),
    .C1(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__o211a_1 _07512_ (.A1(net296),
    .A2(_00413_),
    .B1(_00341_),
    .C1(_00042_),
    .X(_00415_));
 sky130_fd_sc_hd__o21a_1 _07513_ (.A1(_00414_),
    .A2(_00415_),
    .B1(_06402_),
    .X(_00416_));
 sky130_fd_sc_hd__nor3_1 _07514_ (.A(_06402_),
    .B(_00414_),
    .C(_00415_),
    .Y(_00417_));
 sky130_fd_sc_hd__or2_1 _07515_ (.A(_00416_),
    .B(_00417_),
    .X(_00418_));
 sky130_fd_sc_hd__inv_2 _07516_ (.A(_00139_),
    .Y(_00419_));
 sky130_fd_sc_hd__and4b_1 _07517_ (.A_N(_06423_),
    .B(_06425_),
    .C(_03579_),
    .D(_05520_),
    .X(_00420_));
 sky130_fd_sc_hd__buf_2 _07518_ (.A(net81),
    .X(_00421_));
 sky130_fd_sc_hd__a22oi_1 _07519_ (.A1(_03579_),
    .A2(_06410_),
    .B1(_00421_),
    .B2(_02668_),
    .Y(_00422_));
 sky130_fd_sc_hd__and4_1 _07520_ (.A(_03579_),
    .B(_02668_),
    .C(_06410_),
    .D(_00421_),
    .X(_00423_));
 sky130_fd_sc_hd__nor2_1 _07521_ (.A(_00422_),
    .B(_00423_),
    .Y(_00424_));
 sky130_fd_sc_hd__o21a_1 _07522_ (.A1(_06423_),
    .A2(_00420_),
    .B1(_00424_),
    .X(_00425_));
 sky130_fd_sc_hd__nor3_1 _07523_ (.A(_06423_),
    .B(_00420_),
    .C(_00424_),
    .Y(_00426_));
 sky130_fd_sc_hd__nor2_1 _07524_ (.A(_00425_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__and2_1 _07525_ (.A(_06412_),
    .B(_00427_),
    .X(_00428_));
 sky130_fd_sc_hd__nor2_1 _07526_ (.A(_06412_),
    .B(_00427_),
    .Y(_00429_));
 sky130_fd_sc_hd__or2_2 _07527_ (.A(_00428_),
    .B(_00429_),
    .X(_00430_));
 sky130_fd_sc_hd__clkbuf_4 _07528_ (.A(net72),
    .X(_00431_));
 sky130_fd_sc_hd__a22o_1 _07529_ (.A1(_03590_),
    .A2(net71),
    .B1(_00431_),
    .B2(_02657_),
    .X(_00432_));
 sky130_fd_sc_hd__nand4_1 _07530_ (.A(_02657_),
    .B(_03590_),
    .C(_06424_),
    .D(_00431_),
    .Y(_00433_));
 sky130_fd_sc_hd__a22o_1 _07531_ (.A1(_05498_),
    .A2(_05520_),
    .B1(_00432_),
    .B2(_00433_),
    .X(_00434_));
 sky130_fd_sc_hd__nand4_1 _07532_ (.A(_05498_),
    .B(net79),
    .C(_00432_),
    .D(_00433_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_00434_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__inv_2 _07534_ (.A(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__clkbuf_4 _07535_ (.A(net117),
    .X(_00438_));
 sky130_fd_sc_hd__a22o_1 _07536_ (.A1(_05389_),
    .A2(_05444_),
    .B1(_06416_),
    .B2(_03524_),
    .X(_00439_));
 sky130_fd_sc_hd__nand4_2 _07537_ (.A(_03524_),
    .B(_05389_),
    .C(_05444_),
    .D(_06416_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand4_2 _07538_ (.A(_02646_),
    .B(_00438_),
    .C(_00439_),
    .D(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__a22o_1 _07539_ (.A1(_02646_),
    .A2(_00438_),
    .B1(_00439_),
    .B2(_00440_),
    .X(_00442_));
 sky130_fd_sc_hd__nand3_2 _07540_ (.A(_00030_),
    .B(_00441_),
    .C(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__a21o_1 _07541_ (.A1(_00441_),
    .A2(_00442_),
    .B1(_00030_),
    .X(_00444_));
 sky130_fd_sc_hd__and4_1 _07542_ (.A(_03524_),
    .B(_02646_),
    .C(_05444_),
    .D(_06416_),
    .X(_00445_));
 sky130_fd_sc_hd__nor2_1 _07543_ (.A(_00445_),
    .B(_06419_),
    .Y(_00446_));
 sky130_fd_sc_hd__a21oi_1 _07544_ (.A1(_00443_),
    .A2(_00444_),
    .B1(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__a31o_1 _07545_ (.A1(_00443_),
    .A2(_00444_),
    .A3(_00446_),
    .B1(_00447_),
    .X(_00448_));
 sky130_fd_sc_hd__xnor2_2 _07546_ (.A(_00437_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__or2b_1 _07547_ (.A(_06421_),
    .B_N(_06429_),
    .X(_00450_));
 sky130_fd_sc_hd__xor2_2 _07548_ (.A(_00449_),
    .B(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__xor2_2 _07549_ (.A(_00430_),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__clkbuf_4 _07550_ (.A(net177),
    .X(_00453_));
 sky130_fd_sc_hd__clkbuf_4 _07551_ (.A(net107),
    .X(_00454_));
 sky130_fd_sc_hd__a22oi_1 _07552_ (.A1(_03546_),
    .A2(_06437_),
    .B1(_00454_),
    .B2(_02635_),
    .Y(_00455_));
 sky130_fd_sc_hd__and4_1 _07553_ (.A(_02635_),
    .B(_03546_),
    .C(_06437_),
    .D(_00454_),
    .X(_00456_));
 sky130_fd_sc_hd__nor2_1 _07554_ (.A(_00455_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__and3_1 _07555_ (.A(_02745_),
    .B(_00453_),
    .C(_00457_),
    .X(_00458_));
 sky130_fd_sc_hd__a21oi_1 _07556_ (.A1(_02745_),
    .A2(_00453_),
    .B1(_00457_),
    .Y(_00459_));
 sky130_fd_sc_hd__nor2_1 _07557_ (.A(_00458_),
    .B(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _07558_ (.A(net307),
    .B(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__or3_1 _07559_ (.A(_00067_),
    .B(net307),
    .C(_00460_),
    .X(_00462_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(_00067_),
    .B(_00460_),
    .Y(_00463_));
 sky130_fd_sc_hd__and3_1 _07561_ (.A(_00461_),
    .B(_00462_),
    .C(_00463_),
    .X(_00464_));
 sky130_fd_sc_hd__xnor2_1 _07562_ (.A(_00031_),
    .B(_00464_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_00452_),
    .B(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__or2_1 _07564_ (.A(_00452_),
    .B(_00465_),
    .X(_00467_));
 sky130_fd_sc_hd__and3_1 _07565_ (.A(_00075_),
    .B(_00466_),
    .C(_00467_),
    .X(_00468_));
 sky130_fd_sc_hd__a21oi_1 _07566_ (.A1(_00466_),
    .A2(_00467_),
    .B1(_00075_),
    .Y(_00469_));
 sky130_fd_sc_hd__a211oi_2 _07567_ (.A1(_00034_),
    .A2(_00037_),
    .B1(_00468_),
    .C1(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__o211a_1 _07568_ (.A1(_00468_),
    .A2(_00469_),
    .B1(_00034_),
    .C1(_00037_),
    .X(_00471_));
 sky130_fd_sc_hd__a22oi_1 _07569_ (.A1(_05191_),
    .A2(_05202_),
    .B1(_00059_),
    .B2(_03392_),
    .Y(_00472_));
 sky130_fd_sc_hd__and4_1 _07570_ (.A(_03392_),
    .B(_05191_),
    .C(_05202_),
    .D(_00059_),
    .X(_00473_));
 sky130_fd_sc_hd__o2bb2a_1 _07571_ (.A1_N(_03381_),
    .A2_N(_00062_),
    .B1(_00472_),
    .B2(_00473_),
    .X(_00474_));
 sky130_fd_sc_hd__and4bb_1 _07572_ (.A_N(_00472_),
    .B_N(_00473_),
    .C(_03381_),
    .D(_00062_),
    .X(_00475_));
 sky130_fd_sc_hd__a211oi_2 _07573_ (.A1(_00064_),
    .A2(_00066_),
    .B1(_00474_),
    .C1(_00475_),
    .Y(_00476_));
 sky130_fd_sc_hd__o211a_1 _07574_ (.A1(_00474_),
    .A2(_00475_),
    .B1(_00064_),
    .C1(_00066_),
    .X(_00477_));
 sky130_fd_sc_hd__or2_1 _07575_ (.A(_00476_),
    .B(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__clkbuf_4 _07576_ (.A(net123),
    .X(_00479_));
 sky130_fd_sc_hd__clkbuf_4 _07577_ (.A(net195),
    .X(_00480_));
 sky130_fd_sc_hd__buf_2 _07578_ (.A(_00480_),
    .X(_00481_));
 sky130_fd_sc_hd__a22o_1 _07579_ (.A1(_03337_),
    .A2(_00058_),
    .B1(_00481_),
    .B2(net182),
    .X(_00482_));
 sky130_fd_sc_hd__nand4_1 _07580_ (.A(_03337_),
    .B(net182),
    .C(_00058_),
    .D(_00481_),
    .Y(_00483_));
 sky130_fd_sc_hd__and4_1 _07581_ (.A(_02734_),
    .B(_00479_),
    .C(_00482_),
    .D(_00483_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _07582_ (.A1(_02734_),
    .A2(_00479_),
    .B1(_00482_),
    .B2(_00483_),
    .X(_00485_));
 sky130_fd_sc_hd__and2b_1 _07583_ (.A_N(_00484_),
    .B(_00485_),
    .X(_00486_));
 sky130_fd_sc_hd__xnor2_1 _07584_ (.A(_00061_),
    .B(_00486_),
    .Y(_00487_));
 sky130_fd_sc_hd__xor2_1 _07585_ (.A(_00478_),
    .B(_00487_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_2 _07586_ (.A(net186),
    .X(_00489_));
 sky130_fd_sc_hd__a22oi_1 _07587_ (.A1(_03348_),
    .A2(_00049_),
    .B1(_00489_),
    .B2(_02712_),
    .Y(_00490_));
 sky130_fd_sc_hd__and4_1 _07588_ (.A(net191),
    .B(net192),
    .C(_00047_),
    .D(_00489_),
    .X(_00491_));
 sky130_fd_sc_hd__o2bb2a_1 _07589_ (.A1_N(_05115_),
    .A2_N(_05093_),
    .B1(_00490_),
    .B2(_00491_),
    .X(_00492_));
 sky130_fd_sc_hd__and4bb_1 _07590_ (.A_N(_00490_),
    .B_N(_00491_),
    .C(_05115_),
    .D(_05093_),
    .X(_00493_));
 sky130_fd_sc_hd__or2_1 _07591_ (.A(_00492_),
    .B(_00493_),
    .X(_00494_));
 sky130_fd_sc_hd__a41o_1 _07592_ (.A1(_02712_),
    .A2(_03348_),
    .A3(_05115_),
    .A4(_00049_),
    .B1(_00052_),
    .X(_00495_));
 sky130_fd_sc_hd__xnor2_2 _07593_ (.A(_00494_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__a211oi_1 _07594_ (.A1(_05126_),
    .A2(_05147_),
    .B1(_00051_),
    .C1(_00052_),
    .Y(_00497_));
 sky130_fd_sc_hd__or2_1 _07595_ (.A(_00497_),
    .B(_00055_),
    .X(_00498_));
 sky130_fd_sc_hd__xnor2_1 _07596_ (.A(_00496_),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__xnor2_1 _07597_ (.A(_00488_),
    .B(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__xnor2_1 _07598_ (.A(_00093_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__or2_1 _07599_ (.A(_00072_),
    .B(_00501_),
    .X(_00502_));
 sky130_fd_sc_hd__nand2_1 _07600_ (.A(_00072_),
    .B(_00501_),
    .Y(_00503_));
 sky130_fd_sc_hd__and2_1 _07601_ (.A(_00502_),
    .B(_00503_),
    .X(_00504_));
 sky130_fd_sc_hd__inv_2 _07602_ (.A(_00131_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2_1 _07603_ (.A(_04796_),
    .B(_00084_),
    .Y(_00506_));
 sky130_fd_sc_hd__buf_2 _07604_ (.A(net221),
    .X(_00507_));
 sky130_fd_sc_hd__nand4_1 _07605_ (.A(_02855_),
    .B(_03260_),
    .C(_00080_),
    .D(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__nor2_1 _07606_ (.A(_00081_),
    .B(_00508_),
    .Y(_00509_));
 sky130_fd_sc_hd__a22oi_1 _07607_ (.A1(_03260_),
    .A2(_00080_),
    .B1(_00507_),
    .B2(_02855_),
    .Y(_00510_));
 sky130_fd_sc_hd__and2_1 _07608_ (.A(_00081_),
    .B(_00508_),
    .X(_00511_));
 sky130_fd_sc_hd__o32a_1 _07609_ (.A1(_00509_),
    .A2(_00510_),
    .A3(_00511_),
    .B1(_00081_),
    .B2(_04785_),
    .X(_00512_));
 sky130_fd_sc_hd__and4_1 _07610_ (.A(net226),
    .B(_03260_),
    .C(_00080_),
    .D(_00507_),
    .X(_00513_));
 sky130_fd_sc_hd__or4_1 _07611_ (.A(_04785_),
    .B(_00081_),
    .C(_00513_),
    .D(_00510_),
    .X(_00514_));
 sky130_fd_sc_hd__or2b_1 _07612_ (.A(_00512_),
    .B_N(_00514_),
    .X(_00515_));
 sky130_fd_sc_hd__clkbuf_4 _07613_ (.A(net230),
    .X(_00516_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(net217),
    .B(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__and3_1 _07615_ (.A(net218),
    .B(net219),
    .C(net229),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _07616_ (.A1(net219),
    .A2(net228),
    .B1(net229),
    .B2(net218),
    .X(_00519_));
 sky130_fd_sc_hd__a21bo_1 _07617_ (.A1(_04741_),
    .A2(_00518_),
    .B1_N(_00519_),
    .X(_00520_));
 sky130_fd_sc_hd__xor2_1 _07618_ (.A(_00517_),
    .B(_00520_),
    .X(_00521_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(_00088_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__or2_1 _07620_ (.A(_00088_),
    .B(_00521_),
    .X(_00523_));
 sky130_fd_sc_hd__nand2_1 _07621_ (.A(_00522_),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__xor2_1 _07622_ (.A(_00515_),
    .B(_00524_),
    .X(_00525_));
 sky130_fd_sc_hd__o21a_1 _07623_ (.A1(_00506_),
    .A2(_00090_),
    .B1(_00525_),
    .X(_00526_));
 sky130_fd_sc_hd__nor3_1 _07624_ (.A(_00506_),
    .B(_00090_),
    .C(_00525_),
    .Y(_00527_));
 sky130_fd_sc_hd__or2_1 _07625_ (.A(_00526_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__nand3_2 _07626_ (.A(_00106_),
    .B(_00123_),
    .C(_00124_),
    .Y(_00529_));
 sky130_fd_sc_hd__clkbuf_4 _07627_ (.A(net46),
    .X(_00530_));
 sky130_fd_sc_hd__nand2_1 _07628_ (.A(_02822_),
    .B(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(_03084_),
    .B(_00097_),
    .Y(_00532_));
 sky130_fd_sc_hd__and3_1 _07630_ (.A(net42),
    .B(net35),
    .C(net43),
    .X(_00533_));
 sky130_fd_sc_hd__a22o_1 _07631_ (.A1(net35),
    .A2(net43),
    .B1(net36),
    .B2(net42),
    .X(_00534_));
 sky130_fd_sc_hd__a21bo_1 _07632_ (.A1(net36),
    .A2(_00533_),
    .B1_N(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__xor2_1 _07633_ (.A(_00532_),
    .B(_00535_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _07634_ (.A(_00096_),
    .B(_00099_),
    .X(_00537_));
 sky130_fd_sc_hd__xor2_1 _07635_ (.A(_00536_),
    .B(_00537_),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_1 _07636_ (.A(_00531_),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_2 _07637_ (.A(_00103_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__or2_1 _07638_ (.A(_00103_),
    .B(_00539_),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_1 _07639_ (.A(_00540_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__clkbuf_4 _07640_ (.A(net37),
    .X(_00543_));
 sky130_fd_sc_hd__clkbuf_4 _07641_ (.A(net34),
    .X(_00544_));
 sky130_fd_sc_hd__and4_1 _07642_ (.A(_03095_),
    .B(net1),
    .C(_00109_),
    .D(_00544_),
    .X(_00545_));
 sky130_fd_sc_hd__a22oi_1 _07643_ (.A1(_03095_),
    .A2(_00109_),
    .B1(_00544_),
    .B2(_02800_),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_1 _07644_ (.A(_00545_),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__and2_1 _07645_ (.A(net179),
    .B(net12),
    .X(_00548_));
 sky130_fd_sc_hd__buf_6 _07646_ (.A(net190),
    .X(_00549_));
 sky130_fd_sc_hd__buf_6 _07647_ (.A(net201),
    .X(_00550_));
 sky130_fd_sc_hd__nand4_2 _07648_ (.A(_02789_),
    .B(_03106_),
    .C(_00549_),
    .D(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__a22o_1 _07649_ (.A1(net256),
    .A2(net190),
    .B1(net201),
    .B2(net245),
    .X(_00552_));
 sky130_fd_sc_hd__nand3_1 _07650_ (.A(_00548_),
    .B(_00551_),
    .C(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__a21o_1 _07651_ (.A1(_00551_),
    .A2(_00552_),
    .B1(_00548_),
    .X(_00554_));
 sky130_fd_sc_hd__a21bo_1 _07652_ (.A1(_00111_),
    .A2(_00113_),
    .B1_N(_00112_),
    .X(_00555_));
 sky130_fd_sc_hd__nand3_2 _07653_ (.A(_00553_),
    .B(_00554_),
    .C(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__a21o_1 _07654_ (.A1(_00553_),
    .A2(_00554_),
    .B1(_00555_),
    .X(_00557_));
 sky130_fd_sc_hd__nand3_2 _07655_ (.A(_00547_),
    .B(_00556_),
    .C(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__a21o_1 _07656_ (.A1(_00556_),
    .A2(_00557_),
    .B1(_00547_),
    .X(_00559_));
 sky130_fd_sc_hd__o21bai_2 _07657_ (.A1(_00110_),
    .A2(_00118_),
    .B1_N(net315),
    .Y(_00560_));
 sky130_fd_sc_hd__nand3_4 _07658_ (.A(_00558_),
    .B(_00559_),
    .C(_00560_),
    .Y(_00561_));
 sky130_fd_sc_hd__a21o_1 _07659_ (.A1(_00558_),
    .A2(_00559_),
    .B1(_00560_),
    .X(_00562_));
 sky130_fd_sc_hd__nand4_4 _07660_ (.A(_02811_),
    .B(_00543_),
    .C(_00561_),
    .D(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__a22o_1 _07661_ (.A1(_02811_),
    .A2(_00543_),
    .B1(_00561_),
    .B2(_00562_),
    .X(_00564_));
 sky130_fd_sc_hd__and3_1 _07662_ (.A(_00108_),
    .B(_00119_),
    .C(_00120_),
    .X(_00565_));
 sky130_fd_sc_hd__a31o_1 _07663_ (.A1(_02811_),
    .A2(_00107_),
    .A3(_00122_),
    .B1(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__and3_2 _07664_ (.A(_00563_),
    .B(_00564_),
    .C(_00566_),
    .X(_00567_));
 sky130_fd_sc_hd__a21oi_2 _07665_ (.A1(_00563_),
    .A2(_00564_),
    .B1(_00566_),
    .Y(_00568_));
 sky130_fd_sc_hd__nor3_1 _07666_ (.A(_00542_),
    .B(_00567_),
    .C(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__o21a_1 _07667_ (.A1(_00567_),
    .A2(_00568_),
    .B1(_00542_),
    .X(_00570_));
 sky130_fd_sc_hd__a211oi_4 _07668_ (.A1(_00529_),
    .A2(_00127_),
    .B1(net302),
    .C1(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__o211a_1 _07669_ (.A1(_00569_),
    .A2(_00570_),
    .B1(_00529_),
    .C1(_00127_),
    .X(_00572_));
 sky130_fd_sc_hd__nor3_1 _07670_ (.A(_00528_),
    .B(_00571_),
    .C(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__o21a_1 _07671_ (.A1(_00571_),
    .A2(_00572_),
    .B1(_00528_),
    .X(_00574_));
 sky130_fd_sc_hd__a211o_4 _07672_ (.A1(_00505_),
    .A2(_00133_),
    .B1(net299),
    .C1(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__o211ai_4 _07673_ (.A1(net299),
    .A2(_00574_),
    .B1(_00505_),
    .C1(_00133_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand3_4 _07674_ (.A(_00504_),
    .B(_00575_),
    .C(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__a21o_1 _07675_ (.A1(_00575_),
    .A2(_00576_),
    .B1(_00504_),
    .X(_00578_));
 sky130_fd_sc_hd__o211ai_2 _07676_ (.A1(_00135_),
    .A2(net297),
    .B1(_00577_),
    .C1(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__a211o_1 _07677_ (.A1(_00577_),
    .A2(_00578_),
    .B1(_00135_),
    .C1(net297),
    .X(_00580_));
 sky130_fd_sc_hd__or4bb_4 _07678_ (.A(_00470_),
    .B(_00471_),
    .C_N(_00579_),
    .D_N(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__a2bb2o_2 _07679_ (.A1_N(_00470_),
    .A2_N(_00471_),
    .B1(_00579_),
    .B2(_00580_),
    .X(_00582_));
 sky130_fd_sc_hd__o211a_1 _07680_ (.A1(_00419_),
    .A2(_00141_),
    .B1(_00581_),
    .C1(_00582_),
    .X(_00583_));
 sky130_fd_sc_hd__a211oi_4 _07681_ (.A1(_00581_),
    .A2(_00582_),
    .B1(_00419_),
    .C1(_00141_),
    .Y(_00584_));
 sky130_fd_sc_hd__nor3_2 _07682_ (.A(_00418_),
    .B(_00583_),
    .C(net325),
    .Y(_00585_));
 sky130_fd_sc_hd__o21a_1 _07683_ (.A1(_00583_),
    .A2(_00584_),
    .B1(_00418_),
    .X(_00586_));
 sky130_fd_sc_hd__a211o_1 _07684_ (.A1(_00143_),
    .A2(_00145_),
    .B1(_00585_),
    .C1(_00586_),
    .X(_00587_));
 sky130_fd_sc_hd__o211ai_1 _07685_ (.A1(_00585_),
    .A2(_00586_),
    .B1(_00143_),
    .C1(_00145_),
    .Y(_00588_));
 sky130_fd_sc_hd__or4bb_4 _07686_ (.A(_00339_),
    .B(_00340_),
    .C_N(_00587_),
    .D_N(_00588_),
    .X(_00589_));
 sky130_fd_sc_hd__a2bb2o_1 _07687_ (.A1_N(_00339_),
    .A2_N(_00340_),
    .B1(_00587_),
    .B2(_00588_),
    .X(_00590_));
 sky130_fd_sc_hd__o211ai_4 _07688_ (.A1(_00147_),
    .A2(net288),
    .B1(_00589_),
    .C1(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__a211o_1 _07689_ (.A1(_00589_),
    .A2(_00590_),
    .B1(_00147_),
    .C1(net322),
    .X(_00592_));
 sky130_fd_sc_hd__nand3_2 _07690_ (.A(_00192_),
    .B(_00591_),
    .C(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__a21o_1 _07691_ (.A1(_00591_),
    .A2(_00592_),
    .B1(_00192_),
    .X(_00594_));
 sky130_fd_sc_hd__o211ai_4 _07692_ (.A1(_00169_),
    .A2(_00154_),
    .B1(_00593_),
    .C1(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__a211o_1 _07693_ (.A1(_00593_),
    .A2(_00594_),
    .B1(_00169_),
    .C1(_00154_),
    .X(_00596_));
 sky130_fd_sc_hd__o211ai_4 _07694_ (.A1(_06236_),
    .A2(_06240_),
    .B1(_00595_),
    .C1(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__a211o_1 _07695_ (.A1(_00595_),
    .A2(_00596_),
    .B1(_06236_),
    .C1(_06240_),
    .X(_00598_));
 sky130_fd_sc_hd__o211a_1 _07696_ (.A1(_00156_),
    .A2(_00168_),
    .B1(_00597_),
    .C1(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__a211o_1 _07697_ (.A1(_00597_),
    .A2(_00598_),
    .B1(_00156_),
    .C1(_00168_),
    .X(_00600_));
 sky130_fd_sc_hd__or3b_1 _07698_ (.A(_00160_),
    .B(_00599_),
    .C_N(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__o211ai_1 _07699_ (.A1(_00156_),
    .A2(_00168_),
    .B1(_00597_),
    .C1(_00598_),
    .Y(_00602_));
 sky130_fd_sc_hd__and3_1 _07700_ (.A(_06224_),
    .B(_00158_),
    .C(_00159_),
    .X(_00603_));
 sky130_fd_sc_hd__a21o_1 _07701_ (.A1(_00602_),
    .A2(net313),
    .B1(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__and3_1 _07702_ (.A(net280),
    .B(_00601_),
    .C(_00604_),
    .X(_00605_));
 sky130_fd_sc_hd__a21oi_1 _07703_ (.A1(_00601_),
    .A2(_00604_),
    .B1(net280),
    .Y(_00606_));
 sky130_fd_sc_hd__a21boi_1 _07704_ (.A1(_00163_),
    .A2(_00164_),
    .B1_N(_00162_),
    .Y(_00607_));
 sky130_fd_sc_hd__o21ai_1 _07705_ (.A1(_00605_),
    .A2(_00606_),
    .B1(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__or3_1 _07706_ (.A(_00605_),
    .B(_00606_),
    .C(_00607_),
    .X(_00609_));
 sky130_fd_sc_hd__and3_1 _07707_ (.A(_02185_),
    .B(_00608_),
    .C(_00609_),
    .X(_00610_));
 sky130_fd_sc_hd__clkbuf_1 _07708_ (.A(_00610_),
    .X(_00004_));
 sky130_fd_sc_hd__a21oi_1 _07709_ (.A1(_00603_),
    .A2(_00600_),
    .B1(_00599_),
    .Y(_00611_));
 sky130_fd_sc_hd__o21ba_1 _07710_ (.A1(_00170_),
    .A2(_00190_),
    .B1_N(_00189_),
    .X(_00612_));
 sky130_fd_sc_hd__a21oi_2 _07711_ (.A1(_06232_),
    .A2(_00187_),
    .B1(_00185_),
    .Y(_00613_));
 sky130_fd_sc_hd__and4_1 _07712_ (.A(net158),
    .B(net159),
    .C(_06227_),
    .D(_00171_),
    .X(_00614_));
 sky130_fd_sc_hd__a22oi_2 _07713_ (.A1(net159),
    .A2(_06227_),
    .B1(_00171_),
    .B2(_04227_),
    .Y(_00615_));
 sky130_fd_sc_hd__nor2_1 _07714_ (.A(_00614_),
    .B(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__buf_2 _07715_ (.A(net171),
    .X(_00617_));
 sky130_fd_sc_hd__nand2_1 _07716_ (.A(net157),
    .B(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__xnor2_1 _07717_ (.A(_00616_),
    .B(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__or3_1 _07718_ (.A(_00273_),
    .B(_00275_),
    .C(_00619_),
    .X(_00620_));
 sky130_fd_sc_hd__o21a_1 _07719_ (.A1(_00273_),
    .A2(_00275_),
    .B1(_00619_),
    .X(_00621_));
 sky130_fd_sc_hd__inv_2 _07720_ (.A(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(_00620_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _07722_ (.A(_00172_),
    .B(_00175_),
    .Y(_00624_));
 sky130_fd_sc_hd__xnor2_2 _07723_ (.A(_00623_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__xnor2_1 _07724_ (.A(_00178_),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__o21ai_2 _07725_ (.A1(_00281_),
    .A2(_00284_),
    .B1(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__or3_1 _07726_ (.A(_00281_),
    .B(_00284_),
    .C(_00626_),
    .X(_00628_));
 sky130_fd_sc_hd__and2_1 _07727_ (.A(_00627_),
    .B(_00628_),
    .X(_00629_));
 sky130_fd_sc_hd__o21a_1 _07728_ (.A1(_00264_),
    .A2(_00287_),
    .B1(_00629_),
    .X(_00630_));
 sky130_fd_sc_hd__nor3_1 _07729_ (.A(_00264_),
    .B(_00287_),
    .C(_00629_),
    .Y(_00631_));
 sky130_fd_sc_hd__nor2_1 _07730_ (.A(_00630_),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__xor2_1 _07731_ (.A(net303),
    .B(_00632_),
    .X(_00633_));
 sky130_fd_sc_hd__o21a_1 _07732_ (.A1(_00337_),
    .A2(_00339_),
    .B1(_00633_),
    .X(_00634_));
 sky130_fd_sc_hd__nor3_1 _07733_ (.A(_00337_),
    .B(_00339_),
    .C(_00633_),
    .Y(_00635_));
 sky130_fd_sc_hd__nor2_1 _07734_ (.A(_00634_),
    .B(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__xnor2_2 _07735_ (.A(_00613_),
    .B(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__o21ba_1 _07736_ (.A1(_06331_),
    .A2(_00331_),
    .B1_N(_00335_),
    .X(_00638_));
 sky130_fd_sc_hd__nor2_1 _07737_ (.A(_00269_),
    .B(_00276_),
    .Y(_00639_));
 sky130_fd_sc_hd__and2b_1 _07738_ (.A_N(_00268_),
    .B(_00279_),
    .X(_00640_));
 sky130_fd_sc_hd__nor2_1 _07739_ (.A(_06265_),
    .B(_00254_),
    .Y(_00641_));
 sky130_fd_sc_hd__a22o_1 _07740_ (.A1(net166),
    .A2(net161),
    .B1(net162),
    .B2(net165),
    .X(_00642_));
 sky130_fd_sc_hd__inv_2 _07741_ (.A(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__and4_1 _07742_ (.A(_02317_),
    .B(net166),
    .C(net161),
    .D(net162),
    .X(_00644_));
 sky130_fd_sc_hd__o2bb2a_1 _07743_ (.A1_N(net168),
    .A2_N(net160),
    .B1(_00643_),
    .B2(_00644_),
    .X(_00645_));
 sky130_fd_sc_hd__and4b_1 _07744_ (.A_N(_00644_),
    .B(net160),
    .C(net168),
    .D(_00642_),
    .X(_00646_));
 sky130_fd_sc_hd__buf_2 _07745_ (.A(net29),
    .X(_00647_));
 sky130_fd_sc_hd__or4bb_2 _07746_ (.A(_00645_),
    .B(_00646_),
    .C_N(_02207_),
    .D_N(_00647_),
    .X(_00648_));
 sky130_fd_sc_hd__a2bb2o_1 _07747_ (.A1_N(_00645_),
    .A2_N(_00646_),
    .B1(_02207_),
    .B2(_00647_),
    .X(_00649_));
 sky130_fd_sc_hd__and2_1 _07748_ (.A(_00648_),
    .B(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__o21ai_2 _07749_ (.A1(_00252_),
    .A2(_00641_),
    .B1(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__or3_1 _07750_ (.A(_00252_),
    .B(_00641_),
    .C(_00650_),
    .X(_00652_));
 sky130_fd_sc_hd__and2_1 _07751_ (.A(_00651_),
    .B(_00652_),
    .X(_00653_));
 sky130_fd_sc_hd__xnor2_2 _07752_ (.A(_00256_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__xnor2_1 _07753_ (.A(_00278_),
    .B(_00654_),
    .Y(_00655_));
 sky130_fd_sc_hd__xor2_1 _07754_ (.A(_00259_),
    .B(_00655_),
    .X(_00656_));
 sky130_fd_sc_hd__o21ai_1 _07755_ (.A1(_00639_),
    .A2(_00640_),
    .B1(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hd__or3_1 _07756_ (.A(_00639_),
    .B(_00640_),
    .C(_00656_),
    .X(_00658_));
 sky130_fd_sc_hd__nand2_1 _07757_ (.A(_00657_),
    .B(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__or2_1 _07758_ (.A(_00196_),
    .B(_00223_),
    .X(_00660_));
 sky130_fd_sc_hd__nand2_1 _07759_ (.A(_00224_),
    .B(_00262_),
    .Y(_00661_));
 sky130_fd_sc_hd__and2_1 _07760_ (.A(_06323_),
    .B(_00219_),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _07761_ (.A(_00208_),
    .B(_00217_),
    .X(_00663_));
 sky130_fd_sc_hd__or2_1 _07762_ (.A(_00207_),
    .B(_00218_),
    .X(_00664_));
 sky130_fd_sc_hd__buf_2 _07763_ (.A(net136),
    .X(_00665_));
 sky130_fd_sc_hd__a22o_1 _07764_ (.A1(net124),
    .A2(net133),
    .B1(net135),
    .B2(net122),
    .X(_00666_));
 sky130_fd_sc_hd__nand4_2 _07765_ (.A(net122),
    .B(net124),
    .C(net133),
    .D(net135),
    .Y(_00667_));
 sky130_fd_sc_hd__a22o_1 _07766_ (.A1(net121),
    .A2(_00665_),
    .B1(_00666_),
    .B2(_00667_),
    .X(_00668_));
 sky130_fd_sc_hd__nand4_2 _07767_ (.A(net121),
    .B(_00665_),
    .C(_00666_),
    .D(_00667_),
    .Y(_00669_));
 sky130_fd_sc_hd__and3_1 _07768_ (.A(_00203_),
    .B(_00668_),
    .C(_00669_),
    .X(_00670_));
 sky130_fd_sc_hd__a21oi_1 _07769_ (.A1(_00668_),
    .A2(_00669_),
    .B1(_00203_),
    .Y(_00671_));
 sky130_fd_sc_hd__buf_2 _07770_ (.A(net91),
    .X(_00672_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(net94),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__or3_2 _07772_ (.A(_00670_),
    .B(_00671_),
    .C(_00673_),
    .X(_00674_));
 sky130_fd_sc_hd__o21ai_1 _07773_ (.A1(_00670_),
    .A2(_00671_),
    .B1(_00673_),
    .Y(_00675_));
 sky130_fd_sc_hd__and2_1 _07774_ (.A(_00674_),
    .B(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__buf_2 _07775_ (.A(net127),
    .X(_00677_));
 sky130_fd_sc_hd__a22oi_1 _07776_ (.A1(_04314_),
    .A2(_00210_),
    .B1(_00677_),
    .B2(_02218_),
    .Y(_00678_));
 sky130_fd_sc_hd__and4_1 _07777_ (.A(net130),
    .B(net131),
    .C(net126),
    .D(_00677_),
    .X(_00679_));
 sky130_fd_sc_hd__o2bb2a_1 _07778_ (.A1_N(_06151_),
    .A2_N(_06274_),
    .B1(_00678_),
    .B2(_00679_),
    .X(_00680_));
 sky130_fd_sc_hd__and4bb_1 _07779_ (.A_N(_00678_),
    .B_N(_00679_),
    .C(net132),
    .D(_06274_),
    .X(_00681_));
 sky130_fd_sc_hd__nor2_1 _07780_ (.A(_00680_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__a41o_1 _07781_ (.A1(_02218_),
    .A2(_04314_),
    .A3(_06274_),
    .A4(_00210_),
    .B1(_00213_),
    .X(_00683_));
 sky130_fd_sc_hd__xnor2_1 _07782_ (.A(_00682_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__xor2_1 _07783_ (.A(_00215_),
    .B(_00684_),
    .X(_00685_));
 sky130_fd_sc_hd__xnor2_1 _07784_ (.A(_00676_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__xnor2_1 _07785_ (.A(_00323_),
    .B(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__a21o_1 _07786_ (.A1(_00663_),
    .A2(_00664_),
    .B1(_00687_),
    .X(_00688_));
 sky130_fd_sc_hd__nand3_1 _07787_ (.A(_00663_),
    .B(_00664_),
    .C(_00687_),
    .Y(_00689_));
 sky130_fd_sc_hd__o211a_1 _07788_ (.A1(_00662_),
    .A2(_00221_),
    .B1(_00688_),
    .C1(_00689_),
    .X(_00690_));
 sky130_fd_sc_hd__a211oi_1 _07789_ (.A1(_00688_),
    .A2(_00689_),
    .B1(_00662_),
    .C1(_00221_),
    .Y(_00691_));
 sky130_fd_sc_hd__nor2_2 _07790_ (.A(_00690_),
    .B(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__a22o_1 _07791_ (.A1(net26),
    .A2(net18),
    .B1(net27),
    .B2(net17),
    .X(_00693_));
 sky130_fd_sc_hd__nand4_2 _07792_ (.A(_06138_),
    .B(net26),
    .C(net18),
    .D(_06264_),
    .Y(_00694_));
 sky130_fd_sc_hd__a22o_1 _07793_ (.A1(_04435_),
    .A2(net28),
    .B1(_00693_),
    .B2(_00694_),
    .X(_00695_));
 sky130_fd_sc_hd__nand4_1 _07794_ (.A(_04435_),
    .B(_00250_),
    .C(_00693_),
    .D(_00694_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(_00695_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__xnor2_1 _07796_ (.A(_00241_),
    .B(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _07797_ (.A(_00248_),
    .B(_00251_),
    .Y(_00699_));
 sky130_fd_sc_hd__or2b_1 _07798_ (.A(_00698_),
    .B_N(_00699_),
    .X(_00700_));
 sky130_fd_sc_hd__or2b_1 _07799_ (.A(_00699_),
    .B_N(_00698_),
    .X(_00701_));
 sky130_fd_sc_hd__nand2_1 _07800_ (.A(_00700_),
    .B(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__clkbuf_4 _07801_ (.A(net99),
    .X(_00703_));
 sky130_fd_sc_hd__a22o_1 _07802_ (.A1(_04292_),
    .A2(_00238_),
    .B1(_00703_),
    .B2(_02251_),
    .X(_00704_));
 sky130_fd_sc_hd__nand4_2 _07803_ (.A(_04292_),
    .B(net85),
    .C(_00238_),
    .D(_00703_),
    .Y(_00705_));
 sky130_fd_sc_hd__buf_2 _07804_ (.A(net20),
    .X(_00706_));
 sky130_fd_sc_hd__a22o_1 _07805_ (.A1(_04446_),
    .A2(_00239_),
    .B1(_00706_),
    .B2(_02196_),
    .X(_00707_));
 sky130_fd_sc_hd__and4_1 _07806_ (.A(net24),
    .B(net25),
    .C(_00239_),
    .D(_00706_),
    .X(_00708_));
 sky130_fd_sc_hd__inv_2 _07807_ (.A(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__and4_1 _07808_ (.A(_00704_),
    .B(_00705_),
    .C(_00707_),
    .D(_00709_),
    .X(_00710_));
 sky130_fd_sc_hd__a22oi_1 _07809_ (.A1(_00704_),
    .A2(_00705_),
    .B1(_00707_),
    .B2(_00709_),
    .Y(_00711_));
 sky130_fd_sc_hd__or2_1 _07810_ (.A(_00710_),
    .B(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(_00243_),
    .B(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__nor2_1 _07812_ (.A(_00702_),
    .B(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__and2_1 _07813_ (.A(_00702_),
    .B(_00713_),
    .X(_00715_));
 sky130_fd_sc_hd__and2_1 _07814_ (.A(_00231_),
    .B(_00232_),
    .X(_00716_));
 sky130_fd_sc_hd__a22o_1 _07815_ (.A1(net96),
    .A2(net88),
    .B1(net90),
    .B2(net95),
    .X(_00717_));
 sky130_fd_sc_hd__nand4_1 _07816_ (.A(_04413_),
    .B(_06254_),
    .C(net88),
    .D(net90),
    .Y(_00718_));
 sky130_fd_sc_hd__a22oi_1 _07817_ (.A1(_06159_),
    .A2(_06253_),
    .B1(_00717_),
    .B2(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__and4_1 _07818_ (.A(_06159_),
    .B(net97),
    .C(_00717_),
    .D(_00718_),
    .X(_00720_));
 sky130_fd_sc_hd__nor2_1 _07819_ (.A(_00719_),
    .B(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__a41o_1 _07820_ (.A1(_04424_),
    .A2(_06159_),
    .A3(_06134_),
    .A4(_06284_),
    .B1(_00230_),
    .X(_00722_));
 sky130_fd_sc_hd__xnor2_1 _07821_ (.A(_00721_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__nor2_1 _07822_ (.A(_00205_),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__and2_1 _07823_ (.A(_00205_),
    .B(_00723_),
    .X(_00725_));
 sky130_fd_sc_hd__nor2_1 _07824_ (.A(_00724_),
    .B(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__xor2_2 _07825_ (.A(_00716_),
    .B(_00726_),
    .X(_00727_));
 sky130_fd_sc_hd__o21a_1 _07826_ (.A1(_06286_),
    .A2(_00233_),
    .B1(_00235_),
    .X(_00728_));
 sky130_fd_sc_hd__xor2_1 _07827_ (.A(_00727_),
    .B(_00728_),
    .X(_00729_));
 sky130_fd_sc_hd__nor3_1 _07828_ (.A(_00714_),
    .B(_00715_),
    .C(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__o21a_1 _07829_ (.A1(_00714_),
    .A2(_00715_),
    .B1(_00729_),
    .X(_00731_));
 sky130_fd_sc_hd__nor2_1 _07830_ (.A(_00730_),
    .B(_00731_),
    .Y(_00732_));
 sky130_fd_sc_hd__xnor2_2 _07831_ (.A(_00692_),
    .B(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__a21oi_1 _07832_ (.A1(_00660_),
    .A2(_00661_),
    .B1(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__and3_1 _07833_ (.A(_00660_),
    .B(_00661_),
    .C(_00733_),
    .X(_00735_));
 sky130_fd_sc_hd__nor3_1 _07834_ (.A(_00659_),
    .B(_00734_),
    .C(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__o21a_1 _07835_ (.A1(_00734_),
    .A2(_00735_),
    .B1(_00659_),
    .X(_00737_));
 sky130_fd_sc_hd__inv_2 _07836_ (.A(_00383_),
    .Y(_00738_));
 sky130_fd_sc_hd__and2b_1 _07837_ (.A_N(_00290_),
    .B(_00313_),
    .X(_00739_));
 sky130_fd_sc_hd__a21o_1 _07838_ (.A1(_00314_),
    .A2(_00325_),
    .B1(_00739_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_1 _07839_ (.A(_06364_),
    .B(_00347_),
    .Y(_00741_));
 sky130_fd_sc_hd__a22o_1 _07840_ (.A1(net150),
    .A2(net142),
    .B1(net151),
    .B2(net141),
    .X(_00742_));
 sky130_fd_sc_hd__nand4_2 _07841_ (.A(_06177_),
    .B(net150),
    .C(net142),
    .D(net151),
    .Y(_00743_));
 sky130_fd_sc_hd__a22o_1 _07842_ (.A1(net140),
    .A2(net152),
    .B1(_00742_),
    .B2(_00743_),
    .X(_00744_));
 sky130_fd_sc_hd__nand4_1 _07843_ (.A(net140),
    .B(net152),
    .C(_00742_),
    .D(_00743_),
    .Y(_00745_));
 sky130_fd_sc_hd__a21bo_1 _07844_ (.A1(_00316_),
    .A2(_00317_),
    .B1_N(_00315_),
    .X(_00746_));
 sky130_fd_sc_hd__and3_1 _07845_ (.A(_00744_),
    .B(_00745_),
    .C(_00746_),
    .X(_00747_));
 sky130_fd_sc_hd__a21oi_1 _07846_ (.A1(_00744_),
    .A2(_00745_),
    .B1(_00746_),
    .Y(_00748_));
 sky130_fd_sc_hd__clkbuf_4 _07847_ (.A(net153),
    .X(_00749_));
 sky130_fd_sc_hd__a2bb2o_1 _07848_ (.A1_N(_00747_),
    .A2_N(_00748_),
    .B1(_02394_),
    .B2(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__or4bb_1 _07849_ (.A(_00747_),
    .B(_00748_),
    .C_N(net139),
    .D_N(_00749_),
    .X(_00751_));
 sky130_fd_sc_hd__and3_1 _07850_ (.A(_00295_),
    .B(_00750_),
    .C(_00751_),
    .X(_00752_));
 sky130_fd_sc_hd__a21o_1 _07851_ (.A1(_00750_),
    .A2(_00751_),
    .B1(_00295_),
    .X(_00753_));
 sky130_fd_sc_hd__and2b_1 _07852_ (.A_N(_00752_),
    .B(_00753_),
    .X(_00754_));
 sky130_fd_sc_hd__xnor2_2 _07853_ (.A(_00320_),
    .B(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__inv_2 _07854_ (.A(_00310_),
    .Y(_00756_));
 sky130_fd_sc_hd__buf_2 _07855_ (.A(net214),
    .X(_00757_));
 sky130_fd_sc_hd__a22oi_1 _07856_ (.A1(_03941_),
    .A2(_00297_),
    .B1(_00757_),
    .B2(_02459_),
    .Y(_00758_));
 sky130_fd_sc_hd__and4_1 _07857_ (.A(_03941_),
    .B(_02459_),
    .C(_00297_),
    .D(_00757_),
    .X(_00759_));
 sky130_fd_sc_hd__nor2_1 _07858_ (.A(_00758_),
    .B(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__and4_1 _07859_ (.A(_04106_),
    .B(_06077_),
    .C(_06172_),
    .D(_06361_),
    .X(_00761_));
 sky130_fd_sc_hd__and4_1 _07860_ (.A(net200),
    .B(net211),
    .C(_00299_),
    .D(_00300_),
    .X(_00762_));
 sky130_fd_sc_hd__a22o_1 _07861_ (.A1(_06172_),
    .A2(_06361_),
    .B1(net204),
    .B2(net209),
    .X(_00763_));
 sky130_fd_sc_hd__nand4_2 _07862_ (.A(net209),
    .B(_06172_),
    .C(_06361_),
    .D(net204),
    .Y(_00764_));
 sky130_fd_sc_hd__a22o_1 _07863_ (.A1(_06077_),
    .A2(net211),
    .B1(_00763_),
    .B2(_00764_),
    .X(_00765_));
 sky130_fd_sc_hd__nand4_2 _07864_ (.A(_06077_),
    .B(_06304_),
    .C(_00763_),
    .D(_00764_),
    .Y(_00766_));
 sky130_fd_sc_hd__o211ai_2 _07865_ (.A1(_00761_),
    .A2(_00762_),
    .B1(_00765_),
    .C1(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__a211o_1 _07866_ (.A1(_00765_),
    .A2(_00766_),
    .B1(_00761_),
    .C1(_00762_),
    .X(_00768_));
 sky130_fd_sc_hd__nand3_1 _07867_ (.A(_00760_),
    .B(_00767_),
    .C(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21o_1 _07868_ (.A1(_00767_),
    .A2(_00768_),
    .B1(_00760_),
    .X(_00770_));
 sky130_fd_sc_hd__o21bai_1 _07869_ (.A1(_00298_),
    .A2(_00305_),
    .B1_N(_00304_),
    .Y(_00771_));
 sky130_fd_sc_hd__and3_1 _07870_ (.A(_00769_),
    .B(_00770_),
    .C(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__a21oi_1 _07871_ (.A1(_00769_),
    .A2(_00770_),
    .B1(_00771_),
    .Y(_00773_));
 sky130_fd_sc_hd__clkbuf_4 _07872_ (.A(net144),
    .X(_00774_));
 sky130_fd_sc_hd__and4_2 _07873_ (.A(net148),
    .B(net149),
    .C(_00291_),
    .D(_00774_),
    .X(_00775_));
 sky130_fd_sc_hd__and2_1 _07874_ (.A(_00292_),
    .B(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__a22oi_1 _07875_ (.A1(_04139_),
    .A2(_00291_),
    .B1(_00774_),
    .B2(_02383_),
    .Y(_00777_));
 sky130_fd_sc_hd__nor2_2 _07876_ (.A(_00292_),
    .B(_00775_),
    .Y(_00778_));
 sky130_fd_sc_hd__or3_1 _07877_ (.A(_00776_),
    .B(_00777_),
    .C(_00778_),
    .X(_00779_));
 sky130_fd_sc_hd__or3_2 _07878_ (.A(_00772_),
    .B(_00773_),
    .C(_00779_),
    .X(_00780_));
 sky130_fd_sc_hd__o21ai_1 _07879_ (.A1(_00772_),
    .A2(_00773_),
    .B1(_00779_),
    .Y(_00781_));
 sky130_fd_sc_hd__o211a_1 _07880_ (.A1(_00756_),
    .A2(_00311_),
    .B1(_00780_),
    .C1(_00781_),
    .X(_00782_));
 sky130_fd_sc_hd__a211oi_2 _07881_ (.A1(_00780_),
    .A2(_00781_),
    .B1(_00756_),
    .C1(_00311_),
    .Y(_00783_));
 sky130_fd_sc_hd__or3_4 _07882_ (.A(_00755_),
    .B(_00782_),
    .C(_00783_),
    .X(_00784_));
 sky130_fd_sc_hd__o21ai_2 _07883_ (.A1(_00782_),
    .A2(_00783_),
    .B1(_00755_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_2 _07884_ (.A(_00741_),
    .B(_00784_),
    .C(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__a21o_1 _07885_ (.A1(_00784_),
    .A2(_00785_),
    .B1(_00741_),
    .X(_00787_));
 sky130_fd_sc_hd__and3_1 _07886_ (.A(_00740_),
    .B(_00786_),
    .C(_00787_),
    .X(_00788_));
 sky130_fd_sc_hd__a21oi_2 _07887_ (.A1(_00786_),
    .A2(_00787_),
    .B1(_00740_),
    .Y(_00789_));
 sky130_fd_sc_hd__a211oi_4 _07888_ (.A1(_00381_),
    .A2(_00738_),
    .B1(_00788_),
    .C1(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__o211a_1 _07889_ (.A1(_00788_),
    .A2(_00789_),
    .B1(_00381_),
    .C1(_00738_),
    .X(_00791_));
 sky130_fd_sc_hd__nor3_1 _07890_ (.A(_00327_),
    .B(_00790_),
    .C(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__o21a_1 _07891_ (.A1(_00790_),
    .A2(_00791_),
    .B1(_00327_),
    .X(_00793_));
 sky130_fd_sc_hd__nor2_1 _07892_ (.A(_00332_),
    .B(_00330_),
    .Y(_00794_));
 sky130_fd_sc_hd__or4_4 _07893_ (.A(_00329_),
    .B(_00792_),
    .C(_00793_),
    .D(_00794_),
    .X(_00795_));
 sky130_fd_sc_hd__o22ai_4 _07894_ (.A1(net295),
    .A2(_00793_),
    .B1(_00794_),
    .B2(_00329_),
    .Y(_00796_));
 sky130_fd_sc_hd__or4bb_1 _07895_ (.A(net292),
    .B(_00737_),
    .C_N(_00795_),
    .D_N(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__a2bb2o_1 _07896_ (.A1_N(net292),
    .A2_N(_00737_),
    .B1(_00795_),
    .B2(_00796_),
    .X(_00798_));
 sky130_fd_sc_hd__o211a_1 _07897_ (.A1(_00414_),
    .A2(_00417_),
    .B1(_00797_),
    .C1(_00798_),
    .X(_00799_));
 sky130_fd_sc_hd__a211oi_1 _07898_ (.A1(_00797_),
    .A2(_00798_),
    .B1(_00414_),
    .C1(_00417_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor3_1 _07899_ (.A(_00638_),
    .B(_00799_),
    .C(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__o21a_1 _07900_ (.A1(_00799_),
    .A2(_00800_),
    .B1(_00638_),
    .X(_00802_));
 sky130_fd_sc_hd__o211ai_4 _07901_ (.A1(_00419_),
    .A2(_00141_),
    .B1(_00581_),
    .C1(_00582_),
    .Y(_00803_));
 sky130_fd_sc_hd__or3_2 _07902_ (.A(_00418_),
    .B(_00583_),
    .C(net312),
    .X(_00804_));
 sky130_fd_sc_hd__inv_2 _07903_ (.A(_06359_),
    .Y(_00805_));
 sky130_fd_sc_hd__o21ba_1 _07904_ (.A1(_00805_),
    .A2(_00408_),
    .B1_N(_00412_),
    .X(_00806_));
 sky130_fd_sc_hd__inv_2 _07905_ (.A(_00345_),
    .Y(_00807_));
 sky130_fd_sc_hd__nor2_1 _07906_ (.A(_06371_),
    .B(_00377_),
    .Y(_00808_));
 sky130_fd_sc_hd__a32o_1 _07907_ (.A1(_00372_),
    .A2(_00373_),
    .A3(_00375_),
    .B1(_00376_),
    .B2(_00369_),
    .X(_00809_));
 sky130_fd_sc_hd__clkbuf_4 _07908_ (.A(net205),
    .X(_00810_));
 sky130_fd_sc_hd__nand3_2 _07909_ (.A(_02448_),
    .B(_00810_),
    .C(_00368_),
    .Y(_00811_));
 sky130_fd_sc_hd__a21o_1 _07910_ (.A1(_02448_),
    .A2(_00810_),
    .B1(_00368_),
    .X(_00812_));
 sky130_fd_sc_hd__nand2_1 _07911_ (.A(_00811_),
    .B(_00812_),
    .Y(_00813_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(_00809_),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__xnor2_1 _07913_ (.A(_00808_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _07914_ (.A(_00807_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__or2_1 _07915_ (.A(_00807_),
    .B(_00815_),
    .X(_00817_));
 sky130_fd_sc_hd__nand2_1 _07916_ (.A(_00816_),
    .B(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(_06380_),
    .B(_00364_),
    .Y(_00819_));
 sky130_fd_sc_hd__or2_1 _07918_ (.A(_00365_),
    .B(_00378_),
    .X(_00820_));
 sky130_fd_sc_hd__clkbuf_4 _07919_ (.A(net11),
    .X(_00821_));
 sky130_fd_sc_hd__buf_4 _07920_ (.A(net10),
    .X(_00822_));
 sky130_fd_sc_hd__a31o_1 _07921_ (.A1(_02481_),
    .A2(_00822_),
    .A3(_00351_),
    .B1(_00350_),
    .X(_00823_));
 sky130_fd_sc_hd__and3_1 _07922_ (.A(_02481_),
    .B(_00821_),
    .C(_00823_),
    .X(_00824_));
 sky130_fd_sc_hd__a21oi_1 _07923_ (.A1(_02481_),
    .A2(_00821_),
    .B1(_00823_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _07924_ (.A(_00824_),
    .B(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__and3_1 _07925_ (.A(net236),
    .B(net237),
    .C(net248),
    .X(_00827_));
 sky130_fd_sc_hd__a22o_1 _07926_ (.A1(net237),
    .A2(net247),
    .B1(net248),
    .B2(net236),
    .X(_00828_));
 sky130_fd_sc_hd__a21bo_1 _07927_ (.A1(_06383_),
    .A2(_00827_),
    .B1_N(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__clkbuf_4 _07928_ (.A(net249),
    .X(_00830_));
 sky130_fd_sc_hd__nand2_1 _07929_ (.A(_02503_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__xnor2_1 _07930_ (.A(_00829_),
    .B(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__a22o_1 _07931_ (.A1(net244),
    .A2(net239),
    .B1(net240),
    .B2(net243),
    .X(_00833_));
 sky130_fd_sc_hd__clkbuf_4 _07932_ (.A(net239),
    .X(_00834_));
 sky130_fd_sc_hd__nand4_1 _07933_ (.A(_02492_),
    .B(_03864_),
    .C(_00834_),
    .D(net240),
    .Y(_00835_));
 sky130_fd_sc_hd__a22oi_2 _07934_ (.A1(_05969_),
    .A2(_06384_),
    .B1(_00833_),
    .B2(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__and4_2 _07935_ (.A(_05969_),
    .B(_06384_),
    .C(_00833_),
    .D(_00835_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _07936_ (.A(_00836_),
    .B(_00837_),
    .X(_00838_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(_00371_),
    .B(_00372_),
    .Y(_00839_));
 sky130_fd_sc_hd__xnor2_1 _07938_ (.A(_00838_),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__xnor2_1 _07939_ (.A(_00832_),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__and2_1 _07940_ (.A(_00826_),
    .B(_00841_),
    .X(_00842_));
 sky130_fd_sc_hd__nor2_1 _07941_ (.A(_00826_),
    .B(_00841_),
    .Y(_00843_));
 sky130_fd_sc_hd__and2b_1 _07942_ (.A_N(_00363_),
    .B(_00361_),
    .X(_00844_));
 sky130_fd_sc_hd__a22o_1 _07943_ (.A1(net8),
    .A2(net255),
    .B1(net9),
    .B2(net254),
    .X(_00845_));
 sky130_fd_sc_hd__nand4_1 _07944_ (.A(_05914_),
    .B(_05882_),
    .C(_06375_),
    .D(_06368_),
    .Y(_00846_));
 sky130_fd_sc_hd__and2_1 _07945_ (.A(net253),
    .B(net10),
    .X(_00847_));
 sky130_fd_sc_hd__a21o_1 _07946_ (.A1(_00845_),
    .A2(_00846_),
    .B1(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__nand3_1 _07947_ (.A(_00845_),
    .B(_00846_),
    .C(_00847_),
    .Y(_00849_));
 sky130_fd_sc_hd__buf_4 _07948_ (.A(net3),
    .X(_00850_));
 sky130_fd_sc_hd__a22o_1 _07949_ (.A1(_03798_),
    .A2(_00357_),
    .B1(_00850_),
    .B2(_02470_),
    .X(_00851_));
 sky130_fd_sc_hd__and4_2 _07950_ (.A(net6),
    .B(net7),
    .C(net2),
    .D(net3),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_1 _07951_ (.A(_00355_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand4_2 _07952_ (.A(_00848_),
    .B(_00849_),
    .C(_00851_),
    .D(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__a22o_1 _07953_ (.A1(_00848_),
    .A2(_00849_),
    .B1(_00851_),
    .B2(_00853_),
    .X(_00855_));
 sky130_fd_sc_hd__and3_1 _07954_ (.A(_00398_),
    .B(_00854_),
    .C(_00855_),
    .X(_00856_));
 sky130_fd_sc_hd__a21o_1 _07955_ (.A1(_00854_),
    .A2(_00855_),
    .B1(_00398_),
    .X(_00857_));
 sky130_fd_sc_hd__or2b_1 _07956_ (.A(_00856_),
    .B_N(_00857_),
    .X(_00858_));
 sky130_fd_sc_hd__a21bo_1 _07957_ (.A1(_00354_),
    .A2(_00360_),
    .B1_N(_00359_),
    .X(_00859_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(_00858_),
    .B(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__xnor2_1 _07959_ (.A(_00844_),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor3_2 _07960_ (.A(_00842_),
    .B(_00843_),
    .C(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__o21a_1 _07961_ (.A1(_00842_),
    .A2(_00843_),
    .B1(_00861_),
    .X(_00863_));
 sky130_fd_sc_hd__a211oi_2 _07962_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_00862_),
    .C1(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__o211a_1 _07963_ (.A1(_00862_),
    .A2(_00863_),
    .B1(_00819_),
    .C1(_00820_),
    .X(_00865_));
 sky130_fd_sc_hd__nor3_1 _07964_ (.A(_00818_),
    .B(_00864_),
    .C(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__o21a_1 _07965_ (.A1(_00864_),
    .A2(_00865_),
    .B1(_00818_),
    .X(_00867_));
 sky130_fd_sc_hd__or2b_1 _07966_ (.A(_00449_),
    .B_N(_00450_),
    .X(_00868_));
 sky130_fd_sc_hd__o21ai_2 _07967_ (.A1(_00430_),
    .A2(_00451_),
    .B1(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__a32o_1 _07968_ (.A1(_00386_),
    .A2(_00393_),
    .A3(_00394_),
    .B1(_00396_),
    .B2(_00400_),
    .X(_00870_));
 sky130_fd_sc_hd__a21bo_1 _07969_ (.A1(_00388_),
    .A2(_00390_),
    .B1_N(_00389_),
    .X(_00871_));
 sky130_fd_sc_hd__clkbuf_4 _07970_ (.A(net64),
    .X(_00872_));
 sky130_fd_sc_hd__a22oi_1 _07971_ (.A1(_03732_),
    .A2(_00397_),
    .B1(_00872_),
    .B2(net50),
    .Y(_00873_));
 sky130_fd_sc_hd__and4_2 _07972_ (.A(_03732_),
    .B(net50),
    .C(_00397_),
    .D(_00872_),
    .X(_00874_));
 sky130_fd_sc_hd__nor2_1 _07973_ (.A(_00873_),
    .B(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__and2_1 _07974_ (.A(_00871_),
    .B(_00875_),
    .X(_00876_));
 sky130_fd_sc_hd__nor2_1 _07975_ (.A(_00871_),
    .B(_00875_),
    .Y(_00877_));
 sky130_fd_sc_hd__nor2_1 _07976_ (.A(_00876_),
    .B(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__clkbuf_4 _07977_ (.A(net55),
    .X(_00879_));
 sky130_fd_sc_hd__and2_1 _07978_ (.A(net52),
    .B(net62),
    .X(_00880_));
 sky130_fd_sc_hd__a22o_1 _07979_ (.A1(_05761_),
    .A2(net53),
    .B1(_00387_),
    .B2(_03743_),
    .X(_00881_));
 sky130_fd_sc_hd__nand4_2 _07980_ (.A(_03743_),
    .B(_05761_),
    .C(_06343_),
    .D(_00387_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand3_1 _07981_ (.A(_00880_),
    .B(_00881_),
    .C(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hd__a21o_1 _07982_ (.A1(_00881_),
    .A2(_00882_),
    .B1(_00880_),
    .X(_00884_));
 sky130_fd_sc_hd__nand4_2 _07983_ (.A(_02569_),
    .B(_00879_),
    .C(_00883_),
    .D(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__a22o_1 _07984_ (.A1(_02569_),
    .A2(_00879_),
    .B1(_00883_),
    .B2(_00884_),
    .X(_00886_));
 sky130_fd_sc_hd__nand3b_1 _07985_ (.A_N(_00393_),
    .B(_00885_),
    .C(_00886_),
    .Y(_00887_));
 sky130_fd_sc_hd__a21bo_1 _07986_ (.A1(_00885_),
    .A2(_00886_),
    .B1_N(_00393_),
    .X(_00888_));
 sky130_fd_sc_hd__nand3_1 _07987_ (.A(_00878_),
    .B(_00887_),
    .C(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__a21o_1 _07988_ (.A1(_00887_),
    .A2(_00888_),
    .B1(_00878_),
    .X(_00890_));
 sky130_fd_sc_hd__nand3_1 _07989_ (.A(_00428_),
    .B(_00889_),
    .C(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__a21o_1 _07990_ (.A1(_00889_),
    .A2(_00890_),
    .B1(_00428_),
    .X(_00892_));
 sky130_fd_sc_hd__nand3_1 _07991_ (.A(_00870_),
    .B(_00891_),
    .C(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__a21o_1 _07992_ (.A1(_00891_),
    .A2(_00892_),
    .B1(_00870_),
    .X(_00894_));
 sky130_fd_sc_hd__nand2_1 _07993_ (.A(_00893_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__xnor2_1 _07994_ (.A(_00869_),
    .B(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__xnor2_1 _07995_ (.A(_00403_),
    .B(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__a21o_1 _07996_ (.A1(_06357_),
    .A2(_00407_),
    .B1(_00406_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _07997_ (.A(_00897_),
    .B(_00898_),
    .X(_00899_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(_00897_),
    .B(_00898_),
    .Y(_00900_));
 sky130_fd_sc_hd__or4bb_1 _07999_ (.A(net298),
    .B(_00867_),
    .C_N(_00899_),
    .D_N(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__a2bb2o_1 _08000_ (.A1_N(net298),
    .A2_N(_00867_),
    .B1(_00899_),
    .B2(_00900_),
    .X(_00902_));
 sky130_fd_sc_hd__o211a_1 _08001_ (.A1(_00468_),
    .A2(_00470_),
    .B1(_00901_),
    .C1(_00902_),
    .X(_00903_));
 sky130_fd_sc_hd__a211oi_1 _08002_ (.A1(_00901_),
    .A2(_00902_),
    .B1(_00468_),
    .C1(_00470_),
    .Y(_00904_));
 sky130_fd_sc_hd__nor3_2 _08003_ (.A(_00806_),
    .B(_00903_),
    .C(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__o21a_1 _08004_ (.A1(_00903_),
    .A2(_00904_),
    .B1(_00806_),
    .X(_00906_));
 sky130_fd_sc_hd__and2b_1 _08005_ (.A_N(_00031_),
    .B(_00464_),
    .X(_00907_));
 sky130_fd_sc_hd__a21oi_1 _08006_ (.A1(_00452_),
    .A2(_00465_),
    .B1(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand2_1 _08007_ (.A(_00093_),
    .B(_00500_),
    .Y(_00909_));
 sky130_fd_sc_hd__clkbuf_4 _08008_ (.A(net118),
    .X(_00910_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_02646_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__a22o_1 _08010_ (.A1(net77),
    .A2(net72),
    .B1(net73),
    .B2(net76),
    .X(_00912_));
 sky130_fd_sc_hd__nand4_4 _08011_ (.A(_02657_),
    .B(_03590_),
    .C(_00431_),
    .D(net73),
    .Y(_00913_));
 sky130_fd_sc_hd__a22o_1 _08012_ (.A1(_05520_),
    .A2(_06424_),
    .B1(_00912_),
    .B2(_00913_),
    .X(_00914_));
 sky130_fd_sc_hd__nand4_2 _08013_ (.A(net79),
    .B(_06424_),
    .C(_00912_),
    .D(_00913_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_00914_),
    .B(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _08015_ (.A(_00911_),
    .B(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _08016_ (.A(_00911_),
    .B(_00916_),
    .Y(_00918_));
 sky130_fd_sc_hd__and2b_1 _08017_ (.A_N(_00917_),
    .B(_00918_),
    .X(_00919_));
 sky130_fd_sc_hd__nand2_1 _08018_ (.A(_00440_),
    .B(_00441_),
    .Y(_00920_));
 sky130_fd_sc_hd__a22o_1 _08019_ (.A1(_05444_),
    .A2(_06437_),
    .B1(_06416_),
    .B2(_05389_),
    .X(_00921_));
 sky130_fd_sc_hd__nand4_2 _08020_ (.A(_05389_),
    .B(_05444_),
    .C(_06437_),
    .D(_06416_),
    .Y(_00922_));
 sky130_fd_sc_hd__a22o_1 _08021_ (.A1(_03524_),
    .A2(_00438_),
    .B1(_00921_),
    .B2(_00922_),
    .X(_00923_));
 sky130_fd_sc_hd__nand4_2 _08022_ (.A(_03524_),
    .B(_00438_),
    .C(_00921_),
    .D(_00922_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _08023_ (.A(_00456_),
    .B(_00923_),
    .C(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__a21o_1 _08024_ (.A1(_00923_),
    .A2(_00924_),
    .B1(_00456_),
    .X(_00926_));
 sky130_fd_sc_hd__nand3_1 _08025_ (.A(_00920_),
    .B(_00925_),
    .C(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__a21o_1 _08026_ (.A1(_00925_),
    .A2(_00926_),
    .B1(_00920_),
    .X(_00928_));
 sky130_fd_sc_hd__a21bo_1 _08027_ (.A1(_00445_),
    .A2(_00444_),
    .B1_N(_00443_),
    .X(_00929_));
 sky130_fd_sc_hd__nand3_1 _08028_ (.A(_00927_),
    .B(_00928_),
    .C(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__a21o_1 _08029_ (.A1(_00927_),
    .A2(_00928_),
    .B1(_00929_),
    .X(_00931_));
 sky130_fd_sc_hd__nand3_1 _08030_ (.A(_00919_),
    .B(_00930_),
    .C(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__a21o_1 _08031_ (.A1(_00930_),
    .A2(_00931_),
    .B1(_00919_),
    .X(_00933_));
 sky130_fd_sc_hd__a32o_1 _08032_ (.A1(_06419_),
    .A2(_00443_),
    .A3(_00444_),
    .B1(_00448_),
    .B2(_00437_),
    .X(_00934_));
 sky130_fd_sc_hd__nand3_1 _08033_ (.A(_00932_),
    .B(_00933_),
    .C(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__a21o_1 _08034_ (.A1(_00932_),
    .A2(_00933_),
    .B1(_00934_),
    .X(_00936_));
 sky130_fd_sc_hd__clkbuf_4 _08035_ (.A(net82),
    .X(_00937_));
 sky130_fd_sc_hd__a22o_1 _08036_ (.A1(net70),
    .A2(net80),
    .B1(net81),
    .B2(net69),
    .X(_00938_));
 sky130_fd_sc_hd__and4_1 _08037_ (.A(net69),
    .B(net70),
    .C(net80),
    .D(net81),
    .X(_00939_));
 sky130_fd_sc_hd__inv_2 _08038_ (.A(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__a22oi_2 _08039_ (.A1(_02668_),
    .A2(_00937_),
    .B1(_00938_),
    .B2(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__and4b_1 _08040_ (.A_N(_00939_),
    .B(net82),
    .C(net68),
    .D(_00938_),
    .X(_00942_));
 sky130_fd_sc_hd__and2_1 _08041_ (.A(_00433_),
    .B(_00435_),
    .X(_00943_));
 sky130_fd_sc_hd__o21ai_1 _08042_ (.A1(_00941_),
    .A2(_00942_),
    .B1(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__or3_1 _08043_ (.A(_00943_),
    .B(_00941_),
    .C(_00942_),
    .X(_00945_));
 sky130_fd_sc_hd__and2_1 _08044_ (.A(_00944_),
    .B(_00945_),
    .X(_00946_));
 sky130_fd_sc_hd__nor2_1 _08045_ (.A(_00423_),
    .B(_00425_),
    .Y(_00947_));
 sky130_fd_sc_hd__xnor2_2 _08046_ (.A(_00946_),
    .B(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3_1 _08047_ (.A(_00935_),
    .B(_00936_),
    .C(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__a21o_1 _08048_ (.A1(_00935_),
    .A2(_00936_),
    .B1(_00948_),
    .X(_00950_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_00061_),
    .B(_00486_),
    .Y(_00951_));
 sky130_fd_sc_hd__o21ai_1 _08050_ (.A1(_00478_),
    .A2(_00487_),
    .B1(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__clkbuf_4 _08051_ (.A(net178),
    .X(_00953_));
 sky130_fd_sc_hd__a22o_1 _08052_ (.A1(net89),
    .A2(_00453_),
    .B1(_00953_),
    .B2(net78),
    .X(_00954_));
 sky130_fd_sc_hd__nand4_2 _08053_ (.A(_03381_),
    .B(net78),
    .C(_00453_),
    .D(_00953_),
    .Y(_00955_));
 sky130_fd_sc_hd__clkbuf_4 _08054_ (.A(net108),
    .X(_00956_));
 sky130_fd_sc_hd__a22o_1 _08055_ (.A1(net114),
    .A2(_00454_),
    .B1(_00956_),
    .B2(net113),
    .X(_00957_));
 sky130_fd_sc_hd__nand4_2 _08056_ (.A(_02635_),
    .B(_03546_),
    .C(_00454_),
    .D(_00956_),
    .Y(_00958_));
 sky130_fd_sc_hd__and4_1 _08057_ (.A(_00954_),
    .B(_00955_),
    .C(_00957_),
    .D(_00958_),
    .X(_00959_));
 sky130_fd_sc_hd__a22o_1 _08058_ (.A1(_00954_),
    .A2(_00955_),
    .B1(_00957_),
    .B2(_00958_),
    .X(_00960_));
 sky130_fd_sc_hd__or2b_1 _08059_ (.A(_00959_),
    .B_N(_00960_),
    .X(_00961_));
 sky130_fd_sc_hd__xnor2_1 _08060_ (.A(_00476_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__xnor2_1 _08061_ (.A(_00458_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__xor2_1 _08062_ (.A(_00952_),
    .B(_00963_),
    .X(_00964_));
 sky130_fd_sc_hd__xor2_1 _08063_ (.A(_00463_),
    .B(_00964_),
    .X(_00965_));
 sky130_fd_sc_hd__xnor2_1 _08064_ (.A(_00461_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__and3_1 _08065_ (.A(_00949_),
    .B(_00950_),
    .C(_00966_),
    .X(_00967_));
 sky130_fd_sc_hd__a21oi_1 _08066_ (.A1(_00949_),
    .A2(_00950_),
    .B1(_00966_),
    .Y(_00968_));
 sky130_fd_sc_hd__a211oi_2 _08067_ (.A1(_00909_),
    .A2(_00502_),
    .B1(_00967_),
    .C1(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__o211ai_2 _08068_ (.A1(_00967_),
    .A2(_00968_),
    .B1(_00909_),
    .C1(_00502_),
    .Y(_00970_));
 sky130_fd_sc_hd__nor3b_1 _08069_ (.A(_00908_),
    .B(_00969_),
    .C_N(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _08070_ (.A(_00970_),
    .Y(_00972_));
 sky130_fd_sc_hd__o21a_1 _08071_ (.A1(_00969_),
    .A2(_00972_),
    .B1(_00908_),
    .X(_00973_));
 sky130_fd_sc_hd__or2b_1 _08072_ (.A(_00499_),
    .B_N(_00488_),
    .X(_00974_));
 sky130_fd_sc_hd__nand2_1 _08073_ (.A(_00055_),
    .B(_00496_),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_1 _08074_ (.A(_00473_),
    .B(_00475_),
    .Y(_00976_));
 sky130_fd_sc_hd__a22oi_1 _08075_ (.A1(_05202_),
    .A2(_00059_),
    .B1(_00479_),
    .B2(_03392_),
    .Y(_00977_));
 sky130_fd_sc_hd__and4_1 _08076_ (.A(net174),
    .B(net175),
    .C(net111),
    .D(net123),
    .X(_00978_));
 sky130_fd_sc_hd__nor2_1 _08077_ (.A(_00977_),
    .B(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_05191_),
    .B(_00062_),
    .Y(_00980_));
 sky130_fd_sc_hd__xnor2_1 _08079_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__and2b_1 _08080_ (.A_N(_00976_),
    .B(_00981_),
    .X(_00982_));
 sky130_fd_sc_hd__and2b_1 _08081_ (.A_N(_00981_),
    .B(_00976_),
    .X(_00983_));
 sky130_fd_sc_hd__or2_1 _08082_ (.A(_00982_),
    .B(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__clkbuf_4 _08083_ (.A(net134),
    .X(_00985_));
 sky130_fd_sc_hd__nand2_1 _08084_ (.A(_02734_),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__and4_1 _08085_ (.A(net183),
    .B(net182),
    .C(_00058_),
    .D(_00481_),
    .X(_00987_));
 sky130_fd_sc_hd__and2_1 _08086_ (.A(net182),
    .B(net196),
    .X(_00988_));
 sky130_fd_sc_hd__clkbuf_4 _08087_ (.A(net194),
    .X(_00989_));
 sky130_fd_sc_hd__a22o_1 _08088_ (.A1(net184),
    .A2(_00989_),
    .B1(_00480_),
    .B2(net183),
    .X(_00990_));
 sky130_fd_sc_hd__nand4_1 _08089_ (.A(net183),
    .B(net184),
    .C(_00989_),
    .D(_00480_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand3_1 _08090_ (.A(_00988_),
    .B(_00990_),
    .C(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__a21o_1 _08091_ (.A1(_00990_),
    .A2(_00991_),
    .B1(_00988_),
    .X(_00993_));
 sky130_fd_sc_hd__and3_1 _08092_ (.A(_00987_),
    .B(_00992_),
    .C(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__a21oi_1 _08093_ (.A1(_00992_),
    .A2(_00993_),
    .B1(_00987_),
    .Y(_00995_));
 sky130_fd_sc_hd__or3_1 _08094_ (.A(_00986_),
    .B(_00994_),
    .C(_00995_),
    .X(_00996_));
 sky130_fd_sc_hd__o21ai_1 _08095_ (.A1(_00994_),
    .A2(_00995_),
    .B1(_00986_),
    .Y(_00997_));
 sky130_fd_sc_hd__and3_1 _08096_ (.A(_00484_),
    .B(_00996_),
    .C(_00997_),
    .X(_00998_));
 sky130_fd_sc_hd__a21oi_1 _08097_ (.A1(_00996_),
    .A2(_00997_),
    .B1(_00484_),
    .Y(_00999_));
 sky130_fd_sc_hd__nor2_1 _08098_ (.A(_00998_),
    .B(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__xnor2_1 _08099_ (.A(_00984_),
    .B(_01000_),
    .Y(_01001_));
 sky130_fd_sc_hd__buf_2 _08100_ (.A(net187),
    .X(_01002_));
 sky130_fd_sc_hd__a22oi_1 _08101_ (.A1(net192),
    .A2(_00489_),
    .B1(_01002_),
    .B2(net191),
    .Y(_01003_));
 sky130_fd_sc_hd__and4_1 _08102_ (.A(net191),
    .B(net192),
    .C(net186),
    .D(net187),
    .X(_01004_));
 sky130_fd_sc_hd__o2bb2a_1 _08103_ (.A1_N(_05093_),
    .A2_N(_00049_),
    .B1(_01003_),
    .B2(_01004_),
    .X(_01005_));
 sky130_fd_sc_hd__and4bb_1 _08104_ (.A_N(_01003_),
    .B_N(_01004_),
    .C(net193),
    .D(_00049_),
    .X(_01006_));
 sky130_fd_sc_hd__or2_1 _08105_ (.A(_01005_),
    .B(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _08106_ (.A(_00491_),
    .B(_00493_),
    .X(_01008_));
 sky130_fd_sc_hd__xor2_1 _08107_ (.A(_01007_),
    .B(_01008_),
    .X(_01009_));
 sky130_fd_sc_hd__nor2_1 _08108_ (.A(_00522_),
    .B(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _08109_ (.A(_00522_),
    .B(_01009_),
    .Y(_01011_));
 sky130_fd_sc_hd__and2b_1 _08110_ (.A_N(_01010_),
    .B(_01011_),
    .X(_01012_));
 sky130_fd_sc_hd__and2b_1 _08111_ (.A_N(_00494_),
    .B(_00495_),
    .X(_01013_));
 sky130_fd_sc_hd__and2_1 _08112_ (.A(_00497_),
    .B(_00496_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2_1 _08113_ (.A(_01013_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__xnor2_1 _08114_ (.A(_01012_),
    .B(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__xor2_1 _08115_ (.A(_01001_),
    .B(_01016_),
    .X(_01017_));
 sky130_fd_sc_hd__xnor2_1 _08116_ (.A(_00526_),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__a21oi_2 _08117_ (.A1(_00974_),
    .A2(_00975_),
    .B1(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__and3_1 _08118_ (.A(_00974_),
    .B(_00975_),
    .C(_01018_),
    .X(_01020_));
 sky130_fd_sc_hd__o21ai_1 _08119_ (.A1(_00515_),
    .A2(_00524_),
    .B1(_00514_),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _08120_ (.A(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__clkbuf_4 _08121_ (.A(net231),
    .X(_01023_));
 sky130_fd_sc_hd__nand2_1 _08122_ (.A(_02866_),
    .B(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__a22o_1 _08123_ (.A1(net228),
    .A2(net220),
    .B1(net229),
    .B2(net219),
    .X(_01025_));
 sky130_fd_sc_hd__nand4_1 _08124_ (.A(_04752_),
    .B(_04741_),
    .C(net220),
    .D(_00086_),
    .Y(_01026_));
 sky130_fd_sc_hd__nand4_1 _08125_ (.A(_03227_),
    .B(_00516_),
    .C(_01025_),
    .D(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a22o_1 _08126_ (.A1(net218),
    .A2(_00516_),
    .B1(_01025_),
    .B2(_01026_),
    .X(_01028_));
 sky130_fd_sc_hd__a32o_1 _08127_ (.A1(net217),
    .A2(_00516_),
    .A3(_00519_),
    .B1(_00518_),
    .B2(_04741_),
    .X(_01029_));
 sky130_fd_sc_hd__and3_1 _08128_ (.A(_01027_),
    .B(_01028_),
    .C(_01029_),
    .X(_01030_));
 sky130_fd_sc_hd__a21o_1 _08129_ (.A1(_01027_),
    .A2(_01028_),
    .B1(_01029_),
    .X(_01031_));
 sky130_fd_sc_hd__and2b_1 _08130_ (.A_N(_01030_),
    .B(_01031_),
    .X(_01032_));
 sky130_fd_sc_hd__xnor2_1 _08131_ (.A(_01024_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__clkbuf_4 _08132_ (.A(net222),
    .X(_01034_));
 sky130_fd_sc_hd__a22o_1 _08133_ (.A1(_03260_),
    .A2(_00507_),
    .B1(_01034_),
    .B2(_02855_),
    .X(_01035_));
 sky130_fd_sc_hd__nand4_1 _08134_ (.A(_02855_),
    .B(_03260_),
    .C(_00507_),
    .D(_01034_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_1 _08135_ (.A(_00508_),
    .B(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__and4_1 _08136_ (.A(net226),
    .B(_03260_),
    .C(_00507_),
    .D(_01034_),
    .X(_01038_));
 sky130_fd_sc_hd__nand2_1 _08137_ (.A(_00513_),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_1 _08138_ (.A(_01037_),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__and3_1 _08139_ (.A(_00511_),
    .B(_01035_),
    .C(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__a21oi_1 _08140_ (.A1(_01035_),
    .A2(_01040_),
    .B1(_00511_),
    .Y(_01042_));
 sky130_fd_sc_hd__nor2_1 _08141_ (.A(_01041_),
    .B(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__xnor2_1 _08142_ (.A(_01033_),
    .B(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__xnor2_1 _08143_ (.A(_00540_),
    .B(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__xnor2_1 _08144_ (.A(_01022_),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__inv_2 _08145_ (.A(_00567_),
    .Y(_01047_));
 sky130_fd_sc_hd__or3_1 _08146_ (.A(_00542_),
    .B(_00567_),
    .C(_00568_),
    .X(_01048_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(_00536_),
    .B(_00537_),
    .Y(_01049_));
 sky130_fd_sc_hd__or2b_1 _08148_ (.A(_00531_),
    .B_N(_00538_),
    .X(_01050_));
 sky130_fd_sc_hd__buf_4 _08149_ (.A(net47),
    .X(_01051_));
 sky130_fd_sc_hd__a22oi_1 _08150_ (.A1(_03084_),
    .A2(_00530_),
    .B1(_01051_),
    .B2(_02822_),
    .Y(_01052_));
 sky130_fd_sc_hd__and4_1 _08151_ (.A(_03084_),
    .B(net32),
    .C(_00530_),
    .D(_01051_),
    .X(_01053_));
 sky130_fd_sc_hd__nor2_1 _08152_ (.A(_01052_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__and2_1 _08153_ (.A(_04906_),
    .B(_00097_),
    .X(_01055_));
 sky130_fd_sc_hd__a22o_1 _08154_ (.A1(_04862_),
    .A2(net36),
    .B1(net37),
    .B2(_03194_),
    .X(_01056_));
 sky130_fd_sc_hd__nand4_1 _08155_ (.A(_03194_),
    .B(_04862_),
    .C(net36),
    .D(_00543_),
    .Y(_01057_));
 sky130_fd_sc_hd__nand3_1 _08156_ (.A(_01055_),
    .B(_01056_),
    .C(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__a21o_1 _08157_ (.A1(_01056_),
    .A2(_01057_),
    .B1(_01055_),
    .X(_01059_));
 sky130_fd_sc_hd__a32o_1 _08158_ (.A1(_03084_),
    .A2(_00097_),
    .A3(_00534_),
    .B1(_00533_),
    .B2(_00107_),
    .X(_01060_));
 sky130_fd_sc_hd__and3_1 _08159_ (.A(_01058_),
    .B(_01059_),
    .C(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__a21oi_1 _08160_ (.A1(_01058_),
    .A2(_01059_),
    .B1(_01060_),
    .Y(_01062_));
 sky130_fd_sc_hd__nor2_1 _08161_ (.A(_01061_),
    .B(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__xnor2_1 _08162_ (.A(_01054_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_01049_),
    .A2(_01050_),
    .B1(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__inv_2 _08164_ (.A(_01065_),
    .Y(_01066_));
 sky130_fd_sc_hd__and3_1 _08165_ (.A(_01049_),
    .B(_01050_),
    .C(_01064_),
    .X(_01067_));
 sky130_fd_sc_hd__clkbuf_4 _08166_ (.A(net38),
    .X(_01068_));
 sky130_fd_sc_hd__and3_1 _08167_ (.A(net41),
    .B(_01068_),
    .C(_00545_),
    .X(_01069_));
 sky130_fd_sc_hd__a21oi_1 _08168_ (.A1(_02811_),
    .A2(_01068_),
    .B1(_00545_),
    .Y(_01070_));
 sky130_fd_sc_hd__or2_1 _08169_ (.A(_01069_),
    .B(_01070_),
    .X(_01071_));
 sky130_fd_sc_hd__clkbuf_4 _08170_ (.A(net45),
    .X(_01072_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(net1),
    .B(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__and4_1 _08172_ (.A(net112),
    .B(net179),
    .C(net23),
    .D(net34),
    .X(_01074_));
 sky130_fd_sc_hd__a22o_1 _08173_ (.A1(net179),
    .A2(net23),
    .B1(net34),
    .B2(net112),
    .X(_01075_));
 sky130_fd_sc_hd__and2b_1 _08174_ (.A_N(_01074_),
    .B(_01075_),
    .X(_01076_));
 sky130_fd_sc_hd__xnor2_1 _08175_ (.A(_01073_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__and2_1 _08176_ (.A(net12),
    .B(net190),
    .X(_01078_));
 sky130_fd_sc_hd__nand4_1 _08177_ (.A(_02789_),
    .B(_03106_),
    .C(_00550_),
    .D(net212),
    .Y(_01079_));
 sky130_fd_sc_hd__a22o_1 _08178_ (.A1(net256),
    .A2(net201),
    .B1(net212),
    .B2(_02789_),
    .X(_01080_));
 sky130_fd_sc_hd__nand3_1 _08179_ (.A(_01078_),
    .B(_01079_),
    .C(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__a21o_1 _08180_ (.A1(_01079_),
    .A2(_01080_),
    .B1(_01078_),
    .X(_01082_));
 sky130_fd_sc_hd__a21bo_1 _08181_ (.A1(_00548_),
    .A2(_00552_),
    .B1_N(_00551_),
    .X(_01083_));
 sky130_fd_sc_hd__nand3_1 _08182_ (.A(_01081_),
    .B(_01082_),
    .C(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__a21o_1 _08183_ (.A1(_01081_),
    .A2(_01082_),
    .B1(_01083_),
    .X(_01085_));
 sky130_fd_sc_hd__nand3_1 _08184_ (.A(_01077_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__a21o_1 _08185_ (.A1(_01084_),
    .A2(_01085_),
    .B1(_01077_),
    .X(_01087_));
 sky130_fd_sc_hd__a21bo_1 _08186_ (.A1(_00547_),
    .A2(_00557_),
    .B1_N(_00556_),
    .X(_01088_));
 sky130_fd_sc_hd__and3_1 _08187_ (.A(_01086_),
    .B(_01087_),
    .C(_01088_),
    .X(_01089_));
 sky130_fd_sc_hd__a21oi_2 _08188_ (.A1(_01086_),
    .A2(_01087_),
    .B1(_01088_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor3_1 _08189_ (.A(_01071_),
    .B(_01089_),
    .C(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__o21a_1 _08190_ (.A1(_01089_),
    .A2(_01090_),
    .B1(_01071_),
    .X(_01092_));
 sky130_fd_sc_hd__a211oi_4 _08191_ (.A1(_00561_),
    .A2(_00563_),
    .B1(net306),
    .C1(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__o211a_1 _08192_ (.A1(_01091_),
    .A2(_01092_),
    .B1(_00561_),
    .C1(_00563_),
    .X(_01094_));
 sky130_fd_sc_hd__nor4_1 _08193_ (.A(_01066_),
    .B(_01067_),
    .C(_01093_),
    .D(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__o22a_1 _08194_ (.A1(_01066_),
    .A2(_01067_),
    .B1(_01093_),
    .B2(_01094_),
    .X(_01096_));
 sky130_fd_sc_hd__a211oi_2 _08195_ (.A1(_01047_),
    .A2(_01048_),
    .B1(net301),
    .C1(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__o211a_1 _08196_ (.A1(net301),
    .A2(_01096_),
    .B1(_01047_),
    .C1(_01048_),
    .X(_01098_));
 sky130_fd_sc_hd__or3_1 _08197_ (.A(_01046_),
    .B(_01097_),
    .C(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__o21ai_1 _08198_ (.A1(_01097_),
    .A2(_01098_),
    .B1(_01046_),
    .Y(_01100_));
 sky130_fd_sc_hd__o211a_2 _08199_ (.A1(_00571_),
    .A2(net299),
    .B1(_01099_),
    .C1(_01100_),
    .X(_01101_));
 sky130_fd_sc_hd__a211oi_2 _08200_ (.A1(_01099_),
    .A2(_01100_),
    .B1(_00571_),
    .C1(_00573_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor4_1 _08201_ (.A(_01019_),
    .B(_01020_),
    .C(_01101_),
    .D(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__o22a_2 _08202_ (.A1(_01019_),
    .A2(_01020_),
    .B1(_01101_),
    .B2(_01102_),
    .X(_01104_));
 sky130_fd_sc_hd__a211oi_4 _08203_ (.A1(_00575_),
    .A2(_00577_),
    .B1(net294),
    .C1(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__o211a_1 _08204_ (.A1(net294),
    .A2(_01104_),
    .B1(_00575_),
    .C1(_00577_),
    .X(_01106_));
 sky130_fd_sc_hd__nor4_2 _08205_ (.A(_00971_),
    .B(_00973_),
    .C(_01105_),
    .D(_01106_),
    .Y(_01107_));
 sky130_fd_sc_hd__o22a_1 _08206_ (.A1(_00971_),
    .A2(_00973_),
    .B1(_01105_),
    .B2(_01106_),
    .X(_01108_));
 sky130_fd_sc_hd__a211oi_4 _08207_ (.A1(net314),
    .A2(net309),
    .B1(net291),
    .C1(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__o211a_1 _08208_ (.A1(net291),
    .A2(_01108_),
    .B1(net314),
    .C1(net309),
    .X(_01110_));
 sky130_fd_sc_hd__nor4_1 _08209_ (.A(_00905_),
    .B(_00906_),
    .C(_01109_),
    .D(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__o22a_1 _08210_ (.A1(_00905_),
    .A2(_00906_),
    .B1(_01109_),
    .B2(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__a211oi_4 _08211_ (.A1(_00803_),
    .A2(_00804_),
    .B1(net321),
    .C1(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__o211a_1 _08212_ (.A1(net321),
    .A2(_01112_),
    .B1(_00803_),
    .C1(_00804_),
    .X(_01114_));
 sky130_fd_sc_hd__nor4_1 _08213_ (.A(net289),
    .B(_00802_),
    .C(_01113_),
    .D(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__o22a_1 _08214_ (.A1(net289),
    .A2(_00802_),
    .B1(_01113_),
    .B2(_01114_),
    .X(_01116_));
 sky130_fd_sc_hd__a211o_2 _08215_ (.A1(_00587_),
    .A2(_00589_),
    .B1(net287),
    .C1(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__o211ai_2 _08216_ (.A1(net287),
    .A2(_01116_),
    .B1(_00587_),
    .C1(_00589_),
    .Y(_01118_));
 sky130_fd_sc_hd__and3_1 _08217_ (.A(_00637_),
    .B(_01117_),
    .C(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__a21oi_1 _08218_ (.A1(_01117_),
    .A2(_01118_),
    .B1(_00637_),
    .Y(_01120_));
 sky130_fd_sc_hd__a211oi_1 _08219_ (.A1(_00591_),
    .A2(_00593_),
    .B1(_01119_),
    .C1(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__o211a_1 _08220_ (.A1(_01119_),
    .A2(_01120_),
    .B1(_00591_),
    .C1(_00593_),
    .X(_01122_));
 sky130_fd_sc_hd__nor3_1 _08221_ (.A(_00612_),
    .B(_01121_),
    .C(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__o21a_1 _08222_ (.A1(_01121_),
    .A2(_01122_),
    .B1(_00612_),
    .X(_01124_));
 sky130_fd_sc_hd__o211a_1 _08223_ (.A1(_01123_),
    .A2(_01124_),
    .B1(_00595_),
    .C1(_00597_),
    .X(_01125_));
 sky130_fd_sc_hd__a211oi_1 _08224_ (.A1(_00595_),
    .A2(_00597_),
    .B1(_01123_),
    .C1(_01124_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _08225_ (.A(_01125_),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_00611_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__xnor2_1 _08227_ (.A(net281),
    .B(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__o21ba_1 _08228_ (.A1(_00606_),
    .A2(_00607_),
    .B1_N(_00605_),
    .X(_01130_));
 sky130_fd_sc_hd__xnor2_1 _08229_ (.A(_01129_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_00166_),
    .B(_01131_),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _08231_ (.A(_01125_),
    .Y(_01132_));
 sky130_fd_sc_hd__a211o_1 _08232_ (.A1(_00603_),
    .A2(_00600_),
    .B1(_01126_),
    .C1(_00599_),
    .X(_01133_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(_01132_),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__o21bai_1 _08234_ (.A1(_00613_),
    .A2(_00635_),
    .B1_N(_00634_),
    .Y(_01135_));
 sky130_fd_sc_hd__inv_2 _08235_ (.A(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand3_2 _08236_ (.A(_00637_),
    .B(_01117_),
    .C(_01118_),
    .Y(_01137_));
 sky130_fd_sc_hd__a21oi_2 _08237_ (.A1(net303),
    .A2(_00632_),
    .B1(_00630_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_2 _08238_ (.A(_00799_),
    .B(_00801_),
    .Y(_01139_));
 sky130_fd_sc_hd__or2_1 _08239_ (.A(_00734_),
    .B(_00736_),
    .X(_01140_));
 sky130_fd_sc_hd__or2b_1 _08240_ (.A(_00178_),
    .B_N(_00625_),
    .X(_01141_));
 sky130_fd_sc_hd__or2_1 _08241_ (.A(_00259_),
    .B(_00655_),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_1 _08242_ (.A(_00644_),
    .B(_00646_),
    .Y(_01143_));
 sky130_fd_sc_hd__a22oi_1 _08243_ (.A1(net160),
    .A2(net169),
    .B1(_00171_),
    .B2(net159),
    .Y(_01144_));
 sky130_fd_sc_hd__and4_1 _08244_ (.A(net159),
    .B(net160),
    .C(net169),
    .D(net170),
    .X(_01145_));
 sky130_fd_sc_hd__nor2_1 _08245_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__a21oi_1 _08246_ (.A1(_04227_),
    .A2(_00617_),
    .B1(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__and3_1 _08247_ (.A(net158),
    .B(_00617_),
    .C(_01146_),
    .X(_01148_));
 sky130_fd_sc_hd__nor2_1 _08248_ (.A(_01147_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__xnor2_1 _08249_ (.A(_01143_),
    .B(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hd__o21ba_1 _08250_ (.A1(_00615_),
    .A2(_00618_),
    .B1_N(_00614_),
    .X(_01151_));
 sky130_fd_sc_hd__xnor2_1 _08251_ (.A(_01150_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_00172_),
    .B(_00622_),
    .Y(_01153_));
 sky130_fd_sc_hd__and3_1 _08253_ (.A(_00620_),
    .B(_01152_),
    .C(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__a21oi_1 _08254_ (.A1(_00620_),
    .A2(_01153_),
    .B1(_01152_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _08255_ (.A(_01154_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__buf_2 _08256_ (.A(net172),
    .X(_01157_));
 sky130_fd_sc_hd__nand2_1 _08257_ (.A(_02328_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__xnor2_1 _08258_ (.A(_01156_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__nor2_1 _08259_ (.A(_00175_),
    .B(_00623_),
    .Y(_01160_));
 sky130_fd_sc_hd__nand2_2 _08260_ (.A(_01159_),
    .B(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__or2_1 _08261_ (.A(_01159_),
    .B(_01160_),
    .X(_01162_));
 sky130_fd_sc_hd__nand2_1 _08262_ (.A(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__a21oi_1 _08263_ (.A1(_01142_),
    .A2(_00657_),
    .B1(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__and3_1 _08264_ (.A(_01142_),
    .B(_00657_),
    .C(_01163_),
    .X(_01165_));
 sky130_fd_sc_hd__nor2_1 _08265_ (.A(_01164_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__xnor2_2 _08266_ (.A(_01141_),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__xnor2_1 _08267_ (.A(_01140_),
    .B(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_2 _08268_ (.A(_00627_),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__and2_1 _08269_ (.A(_00627_),
    .B(_01168_),
    .X(_01170_));
 sky130_fd_sc_hd__nor2_1 _08270_ (.A(_01169_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__xnor2_2 _08271_ (.A(_01139_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__xnor2_2 _08272_ (.A(_01138_),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _08273_ (.A(_00795_),
    .B(_00797_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _08274_ (.A(_00256_),
    .B(_00653_),
    .Y(_01175_));
 sky130_fd_sc_hd__o21ai_2 _08275_ (.A1(_00278_),
    .A2(_00654_),
    .B1(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__and2b_1 _08276_ (.A_N(_00728_),
    .B(_00727_),
    .X(_01177_));
 sky130_fd_sc_hd__or2_1 _08277_ (.A(_01177_),
    .B(_00730_),
    .X(_01178_));
 sky130_fd_sc_hd__o21bai_2 _08278_ (.A1(_00243_),
    .A2(_00712_),
    .B1_N(_00714_),
    .Y(_01179_));
 sky130_fd_sc_hd__or2_1 _08279_ (.A(_00241_),
    .B(_00697_),
    .X(_01180_));
 sky130_fd_sc_hd__buf_2 _08280_ (.A(net30),
    .X(_01181_));
 sky130_fd_sc_hd__a22o_1 _08281_ (.A1(_04435_),
    .A2(_00647_),
    .B1(_01181_),
    .B2(net15),
    .X(_01182_));
 sky130_fd_sc_hd__and4_1 _08282_ (.A(net16),
    .B(net15),
    .C(net29),
    .D(_01181_),
    .X(_01183_));
 sky130_fd_sc_hd__inv_2 _08283_ (.A(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__and2_1 _08284_ (.A(_01182_),
    .B(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__a22o_1 _08285_ (.A1(net166),
    .A2(net162),
    .B1(net163),
    .B2(net165),
    .X(_01186_));
 sky130_fd_sc_hd__inv_2 _08286_ (.A(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__buf_2 _08287_ (.A(net163),
    .X(_01188_));
 sky130_fd_sc_hd__and4_1 _08288_ (.A(_02317_),
    .B(_04238_),
    .C(net162),
    .D(_01188_),
    .X(_01189_));
 sky130_fd_sc_hd__o2bb2a_1 _08289_ (.A1_N(net168),
    .A2_N(_00270_),
    .B1(_01187_),
    .B2(_01189_),
    .X(_01190_));
 sky130_fd_sc_hd__and4b_1 _08290_ (.A_N(_01189_),
    .B(_00270_),
    .C(net168),
    .D(_01186_),
    .X(_01191_));
 sky130_fd_sc_hd__nor2_1 _08291_ (.A(_01190_),
    .B(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__xnor2_1 _08292_ (.A(_01185_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__a21oi_1 _08293_ (.A1(_01180_),
    .A2(_00700_),
    .B1(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__and3_1 _08294_ (.A(_01180_),
    .B(_00700_),
    .C(_01193_),
    .X(_01195_));
 sky130_fd_sc_hd__or2_1 _08295_ (.A(_01194_),
    .B(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__xor2_2 _08296_ (.A(_00648_),
    .B(_01196_),
    .X(_01197_));
 sky130_fd_sc_hd__xnor2_2 _08297_ (.A(_01179_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__xor2_2 _08298_ (.A(_00651_),
    .B(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__xnor2_2 _08299_ (.A(_01178_),
    .B(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__xor2_2 _08300_ (.A(_01176_),
    .B(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__a22o_1 _08301_ (.A1(_06261_),
    .A2(_06264_),
    .B1(net19),
    .B2(_06142_),
    .X(_01202_));
 sky130_fd_sc_hd__nand4_2 _08302_ (.A(_06142_),
    .B(_06261_),
    .C(_06264_),
    .D(_00239_),
    .Y(_01203_));
 sky130_fd_sc_hd__a22o_1 _08303_ (.A1(_06138_),
    .A2(_00250_),
    .B1(_01202_),
    .B2(_01203_),
    .X(_01204_));
 sky130_fd_sc_hd__nand4_1 _08304_ (.A(_06138_),
    .B(_00250_),
    .C(_01202_),
    .D(_01203_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _08305_ (.A(_01204_),
    .B(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_00709_),
    .B(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__a21oi_1 _08307_ (.A1(_00694_),
    .A2(_00696_),
    .B1(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__and3_1 _08308_ (.A(_00694_),
    .B(_00696_),
    .C(_01207_),
    .X(_01209_));
 sky130_fd_sc_hd__or2_1 _08309_ (.A(_01208_),
    .B(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__a22oi_1 _08310_ (.A1(net87),
    .A2(net98),
    .B1(net99),
    .B2(net86),
    .Y(_01211_));
 sky130_fd_sc_hd__and4_1 _08311_ (.A(net86),
    .B(net87),
    .C(net98),
    .D(net99),
    .X(_01212_));
 sky130_fd_sc_hd__o2bb2a_1 _08312_ (.A1_N(net85),
    .A2_N(net101),
    .B1(_01211_),
    .B2(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__and4bb_1 _08313_ (.A_N(_01211_),
    .B_N(_01212_),
    .C(net85),
    .D(net101),
    .X(_01214_));
 sky130_fd_sc_hd__or2_1 _08314_ (.A(_01213_),
    .B(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_1 _08315_ (.A(_00705_),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__buf_2 _08316_ (.A(net21),
    .X(_01217_));
 sky130_fd_sc_hd__a22o_1 _08317_ (.A1(_04446_),
    .A2(_00706_),
    .B1(_01217_),
    .B2(_02196_),
    .X(_01218_));
 sky130_fd_sc_hd__inv_2 _08318_ (.A(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__and4_1 _08319_ (.A(_02196_),
    .B(_04446_),
    .C(_00706_),
    .D(_01217_),
    .X(_01220_));
 sky130_fd_sc_hd__nor2_1 _08320_ (.A(_01219_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__xnor2_1 _08321_ (.A(_01216_),
    .B(_01221_),
    .Y(_01222_));
 sky130_fd_sc_hd__xnor2_1 _08322_ (.A(_00710_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__or2_1 _08323_ (.A(_01210_),
    .B(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(_01210_),
    .B(_01223_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_01224_),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__and2_1 _08326_ (.A(_00721_),
    .B(_00722_),
    .X(_01227_));
 sky130_fd_sc_hd__nand3_1 _08327_ (.A(_00203_),
    .B(_00668_),
    .C(_00669_),
    .Y(_01228_));
 sky130_fd_sc_hd__and4_1 _08328_ (.A(_04424_),
    .B(_06134_),
    .C(_06284_),
    .D(_00200_),
    .X(_01229_));
 sky130_fd_sc_hd__a22o_1 _08329_ (.A1(_06254_),
    .A2(net90),
    .B1(net91),
    .B2(_04413_),
    .X(_01230_));
 sky130_fd_sc_hd__nand4_2 _08330_ (.A(_04413_),
    .B(_06254_),
    .C(net90),
    .D(net91),
    .Y(_01231_));
 sky130_fd_sc_hd__a22o_1 _08331_ (.A1(_06284_),
    .A2(net97),
    .B1(_01230_),
    .B2(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__nand4_2 _08332_ (.A(_06284_),
    .B(_06253_),
    .C(_01230_),
    .D(_01231_),
    .Y(_01233_));
 sky130_fd_sc_hd__o211a_1 _08333_ (.A1(_01229_),
    .A2(_00720_),
    .B1(_01232_),
    .C1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__a211oi_1 _08334_ (.A1(_01232_),
    .A2(_01233_),
    .B1(_01229_),
    .C1(_00720_),
    .Y(_01235_));
 sky130_fd_sc_hd__or2_1 _08335_ (.A(_01234_),
    .B(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__a21oi_2 _08336_ (.A1(_01228_),
    .A2(_00674_),
    .B1(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__and3_1 _08337_ (.A(_01228_),
    .B(_00674_),
    .C(_01236_),
    .X(_01238_));
 sky130_fd_sc_hd__nor2_1 _08338_ (.A(_01237_),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__xnor2_2 _08339_ (.A(_01227_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__a21oi_2 _08340_ (.A1(_00716_),
    .A2(_00726_),
    .B1(_00724_),
    .Y(_01241_));
 sky130_fd_sc_hd__xnor2_1 _08341_ (.A(_01240_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _08342_ (.A(_01226_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__and2_1 _08343_ (.A(_01226_),
    .B(_01242_),
    .X(_01244_));
 sky130_fd_sc_hd__or2_2 _08344_ (.A(_01243_),
    .B(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__or2_1 _08345_ (.A(_00323_),
    .B(_00686_),
    .X(_01246_));
 sky130_fd_sc_hd__nor2_1 _08346_ (.A(_00215_),
    .B(_00684_),
    .Y(_01247_));
 sky130_fd_sc_hd__a21o_1 _08347_ (.A1(_00676_),
    .A2(_00685_),
    .B1(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__a21oi_2 _08348_ (.A1(_00320_),
    .A2(_00753_),
    .B1(_00752_),
    .Y(_01249_));
 sky130_fd_sc_hd__buf_2 _08349_ (.A(net137),
    .X(_01250_));
 sky130_fd_sc_hd__clkbuf_4 _08350_ (.A(net92),
    .X(_01251_));
 sky130_fd_sc_hd__a22oi_2 _08351_ (.A1(_02229_),
    .A2(_01250_),
    .B1(_01251_),
    .B2(net94),
    .Y(_01252_));
 sky130_fd_sc_hd__and4_2 _08352_ (.A(net121),
    .B(net94),
    .C(_01250_),
    .D(_01251_),
    .X(_01253_));
 sky130_fd_sc_hd__nor2_1 _08353_ (.A(_01252_),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__a22o_1 _08354_ (.A1(net125),
    .A2(_06283_),
    .B1(_00201_),
    .B2(net124),
    .X(_01255_));
 sky130_fd_sc_hd__nand4_1 _08355_ (.A(net124),
    .B(net125),
    .C(_06283_),
    .D(_00201_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _08356_ (.A(_01255_),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__and2_1 _08357_ (.A(_04303_),
    .B(_00665_),
    .X(_01258_));
 sky130_fd_sc_hd__xor2_1 _08358_ (.A(_01257_),
    .B(_01258_),
    .X(_01259_));
 sky130_fd_sc_hd__nand2_1 _08359_ (.A(_00667_),
    .B(_00669_),
    .Y(_01260_));
 sky130_fd_sc_hd__xor2_1 _08360_ (.A(_01259_),
    .B(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__xor2_1 _08361_ (.A(_01254_),
    .B(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__nand2_1 _08362_ (.A(_00682_),
    .B(_00683_),
    .Y(_01263_));
 sky130_fd_sc_hd__clkbuf_4 _08363_ (.A(net128),
    .X(_01264_));
 sky130_fd_sc_hd__and3_1 _08364_ (.A(net130),
    .B(net131),
    .C(net127),
    .X(_01265_));
 sky130_fd_sc_hd__a22o_1 _08365_ (.A1(net131),
    .A2(net127),
    .B1(net128),
    .B2(net130),
    .X(_01266_));
 sky130_fd_sc_hd__a21bo_1 _08366_ (.A1(_01264_),
    .A2(_01265_),
    .B1_N(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__nand2_1 _08367_ (.A(_06151_),
    .B(_00210_),
    .Y(_01268_));
 sky130_fd_sc_hd__xor2_1 _08368_ (.A(_01267_),
    .B(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__nor2_1 _08369_ (.A(_00679_),
    .B(_00681_),
    .Y(_01270_));
 sky130_fd_sc_hd__xor2_1 _08370_ (.A(_01269_),
    .B(_01270_),
    .X(_01271_));
 sky130_fd_sc_hd__xnor2_1 _08371_ (.A(_01263_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__xnor2_1 _08372_ (.A(_01262_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__xnor2_1 _08373_ (.A(_01249_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__xor2_1 _08374_ (.A(_01248_),
    .B(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__a21oi_2 _08375_ (.A1(_01246_),
    .A2(_00688_),
    .B1(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__and3_1 _08376_ (.A(_01246_),
    .B(_00688_),
    .C(_01275_),
    .X(_01277_));
 sky130_fd_sc_hd__or2_2 _08377_ (.A(_01276_),
    .B(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__xnor2_4 _08378_ (.A(_01245_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__a21o_1 _08379_ (.A1(_00692_),
    .A2(_00732_),
    .B1(_00690_),
    .X(_01280_));
 sky130_fd_sc_hd__xor2_2 _08380_ (.A(_01279_),
    .B(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__xnor2_2 _08381_ (.A(_01201_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__inv_2 _08382_ (.A(_00786_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _08383_ (.A(_01283_),
    .B(_00788_),
    .Y(_01284_));
 sky130_fd_sc_hd__inv_2 _08384_ (.A(_00782_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_1 _08385_ (.A(_00808_),
    .B(_00814_),
    .Y(_01286_));
 sky130_fd_sc_hd__or2b_1 _08386_ (.A(_00747_),
    .B_N(_00751_),
    .X(_01287_));
 sky130_fd_sc_hd__buf_2 _08387_ (.A(net154),
    .X(_01288_));
 sky130_fd_sc_hd__a22oi_1 _08388_ (.A1(_04128_),
    .A2(_00749_),
    .B1(_01288_),
    .B2(_02394_),
    .Y(_01289_));
 sky130_fd_sc_hd__and4_1 _08389_ (.A(_04128_),
    .B(net139),
    .C(_00749_),
    .D(_01288_),
    .X(_01290_));
 sky130_fd_sc_hd__nor2_1 _08390_ (.A(_01289_),
    .B(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__and4_1 _08391_ (.A(_06178_),
    .B(_06171_),
    .C(_06311_),
    .D(_06319_),
    .X(_01292_));
 sky130_fd_sc_hd__clkbuf_4 _08392_ (.A(net152),
    .X(_01293_));
 sky130_fd_sc_hd__and4_1 _08393_ (.A(_04128_),
    .B(_01293_),
    .C(_00742_),
    .D(_00743_),
    .X(_01294_));
 sky130_fd_sc_hd__a22o_1 _08394_ (.A1(net142),
    .A2(_06319_),
    .B1(_00291_),
    .B2(_06171_),
    .X(_01295_));
 sky130_fd_sc_hd__nand4_4 _08395_ (.A(_06171_),
    .B(_06311_),
    .C(_06319_),
    .D(_00291_),
    .Y(_01296_));
 sky130_fd_sc_hd__a22o_1 _08396_ (.A1(_06178_),
    .A2(_01293_),
    .B1(_01295_),
    .B2(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__nand4_4 _08397_ (.A(_06177_),
    .B(_01293_),
    .C(_01295_),
    .D(_01296_),
    .Y(_01298_));
 sky130_fd_sc_hd__o211ai_2 _08398_ (.A1(_01292_),
    .A2(_01294_),
    .B1(_01297_),
    .C1(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__a211o_1 _08399_ (.A1(_01297_),
    .A2(_01298_),
    .B1(_01292_),
    .C1(_01294_),
    .X(_01300_));
 sky130_fd_sc_hd__nand3_2 _08400_ (.A(_01291_),
    .B(_01299_),
    .C(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__a21o_1 _08401_ (.A1(_01299_),
    .A2(_01300_),
    .B1(_01291_),
    .X(_01302_));
 sky130_fd_sc_hd__nand3_4 _08402_ (.A(_00778_),
    .B(_01301_),
    .C(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__a21o_1 _08403_ (.A1(_01301_),
    .A2(_01302_),
    .B1(_00778_),
    .X(_01304_));
 sky130_fd_sc_hd__nand3_4 _08404_ (.A(_01287_),
    .B(_01303_),
    .C(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__a21o_1 _08405_ (.A1(_01303_),
    .A2(_01304_),
    .B1(_01287_),
    .X(_01306_));
 sky130_fd_sc_hd__nand2_2 _08406_ (.A(_01305_),
    .B(_01306_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand3_1 _08407_ (.A(_00769_),
    .B(_00770_),
    .C(_00771_),
    .Y(_01308_));
 sky130_fd_sc_hd__clkbuf_4 _08408_ (.A(net146),
    .X(_01309_));
 sky130_fd_sc_hd__a22o_1 _08409_ (.A1(net149),
    .A2(_00774_),
    .B1(_01309_),
    .B2(_02383_),
    .X(_01310_));
 sky130_fd_sc_hd__and4_1 _08410_ (.A(net148),
    .B(net149),
    .C(net144),
    .D(net146),
    .X(_01311_));
 sky130_fd_sc_hd__inv_2 _08411_ (.A(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__and3_1 _08412_ (.A(_00759_),
    .B(_01310_),
    .C(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__a21o_1 _08413_ (.A1(_01310_),
    .A2(_01312_),
    .B1(_00759_),
    .X(_01314_));
 sky130_fd_sc_hd__or2b_1 _08414_ (.A(_01313_),
    .B_N(_01314_),
    .X(_01315_));
 sky130_fd_sc_hd__xor2_2 _08415_ (.A(_00775_),
    .B(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__a22oi_2 _08416_ (.A1(_06077_),
    .A2(net213),
    .B1(net214),
    .B2(_03941_),
    .Y(_01317_));
 sky130_fd_sc_hd__and4_1 _08417_ (.A(net200),
    .B(_06077_),
    .C(net213),
    .D(net214),
    .X(_01318_));
 sky130_fd_sc_hd__nor2_1 _08418_ (.A(_01317_),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_1 _08419_ (.A(_02459_),
    .B(net215),
    .Y(_01320_));
 sky130_fd_sc_hd__xnor2_1 _08420_ (.A(_01319_),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__and4_1 _08421_ (.A(_04106_),
    .B(_06173_),
    .C(_06362_),
    .D(_00343_),
    .X(_01322_));
 sky130_fd_sc_hd__and4_1 _08422_ (.A(_06086_),
    .B(_06304_),
    .C(_00763_),
    .D(_00764_),
    .X(_01323_));
 sky130_fd_sc_hd__a22o_1 _08423_ (.A1(_06172_),
    .A2(net204),
    .B1(net205),
    .B2(net209),
    .X(_01324_));
 sky130_fd_sc_hd__nand4_1 _08424_ (.A(_04106_),
    .B(_06172_),
    .C(net204),
    .D(net205),
    .Y(_01325_));
 sky130_fd_sc_hd__a22o_1 _08425_ (.A1(_06362_),
    .A2(_06304_),
    .B1(_01324_),
    .B2(_01325_),
    .X(_01326_));
 sky130_fd_sc_hd__nand4_1 _08426_ (.A(_06362_),
    .B(_06304_),
    .C(_01324_),
    .D(_01325_),
    .Y(_01327_));
 sky130_fd_sc_hd__o211ai_2 _08427_ (.A1(_01322_),
    .A2(_01323_),
    .B1(_01326_),
    .C1(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hd__a211o_1 _08428_ (.A1(_01326_),
    .A2(_01327_),
    .B1(_01322_),
    .C1(_01323_),
    .X(_01329_));
 sky130_fd_sc_hd__nand3_1 _08429_ (.A(_01321_),
    .B(_01328_),
    .C(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__a21o_1 _08430_ (.A1(_01328_),
    .A2(_01329_),
    .B1(_01321_),
    .X(_01331_));
 sky130_fd_sc_hd__a21bo_1 _08431_ (.A1(_00760_),
    .A2(_00768_),
    .B1_N(_00767_),
    .X(_01332_));
 sky130_fd_sc_hd__and3_1 _08432_ (.A(_01330_),
    .B(_01331_),
    .C(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__a21oi_1 _08433_ (.A1(_01330_),
    .A2(_01331_),
    .B1(_01332_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor3_2 _08434_ (.A(_01316_),
    .B(_01333_),
    .C(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__o21a_1 _08435_ (.A1(_01333_),
    .A2(_01334_),
    .B1(_01316_),
    .X(_01336_));
 sky130_fd_sc_hd__a211oi_2 _08436_ (.A1(_01308_),
    .A2(_00780_),
    .B1(_01335_),
    .C1(_01336_),
    .Y(_01337_));
 sky130_fd_sc_hd__o211a_1 _08437_ (.A1(_01335_),
    .A2(_01336_),
    .B1(_01308_),
    .C1(_00780_),
    .X(_01338_));
 sky130_fd_sc_hd__nor3_2 _08438_ (.A(_01307_),
    .B(_01337_),
    .C(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__o21a_1 _08439_ (.A1(_01337_),
    .A2(_01338_),
    .B1(_01307_),
    .X(_01340_));
 sky130_fd_sc_hd__a211oi_2 _08440_ (.A1(_01286_),
    .A2(_00817_),
    .B1(_01339_),
    .C1(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o211a_1 _08441_ (.A1(_01339_),
    .A2(_01340_),
    .B1(_01286_),
    .C1(_00817_),
    .X(_01342_));
 sky130_fd_sc_hd__a211o_1 _08442_ (.A1(_01285_),
    .A2(_00784_),
    .B1(_01341_),
    .C1(_01342_),
    .X(_01343_));
 sky130_fd_sc_hd__o211ai_2 _08443_ (.A1(_01341_),
    .A2(_01342_),
    .B1(_01285_),
    .C1(_00784_),
    .Y(_01344_));
 sky130_fd_sc_hd__o211a_2 _08444_ (.A1(_00864_),
    .A2(_00866_),
    .B1(_01343_),
    .C1(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__a211oi_2 _08445_ (.A1(_01343_),
    .A2(_01344_),
    .B1(_00864_),
    .C1(_00866_),
    .Y(_01346_));
 sky130_fd_sc_hd__or3_1 _08446_ (.A(_01284_),
    .B(_01345_),
    .C(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__o21ai_1 _08447_ (.A1(_01345_),
    .A2(_01346_),
    .B1(_01284_),
    .Y(_01348_));
 sky130_fd_sc_hd__o211a_1 _08448_ (.A1(_00790_),
    .A2(net295),
    .B1(_01347_),
    .C1(_01348_),
    .X(_01349_));
 sky130_fd_sc_hd__a211oi_2 _08449_ (.A1(_01347_),
    .A2(_01348_),
    .B1(_00790_),
    .C1(net295),
    .Y(_01350_));
 sky130_fd_sc_hd__or3_1 _08450_ (.A(_01282_),
    .B(_01349_),
    .C(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__o21ai_1 _08451_ (.A1(_01349_),
    .A2(_01350_),
    .B1(_01282_),
    .Y(_01352_));
 sky130_fd_sc_hd__o211ai_2 _08452_ (.A1(_00903_),
    .A2(_00905_),
    .B1(_01351_),
    .C1(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__a211o_1 _08453_ (.A1(_01351_),
    .A2(_01352_),
    .B1(_00903_),
    .C1(_00905_),
    .X(_01354_));
 sky130_fd_sc_hd__nand3_1 _08454_ (.A(_01174_),
    .B(_01353_),
    .C(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__a21o_1 _08455_ (.A1(_01353_),
    .A2(_01354_),
    .B1(_01174_),
    .X(_01356_));
 sky130_fd_sc_hd__nand2_1 _08456_ (.A(_00899_),
    .B(_00901_),
    .Y(_01357_));
 sky130_fd_sc_hd__or2_2 _08457_ (.A(_00969_),
    .B(_00971_),
    .X(_01358_));
 sky130_fd_sc_hd__and3_1 _08458_ (.A(_00809_),
    .B(_00811_),
    .C(_00812_),
    .X(_01359_));
 sky130_fd_sc_hd__inv_2 _08459_ (.A(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__o211a_1 _08460_ (.A1(_00836_),
    .A2(_00837_),
    .B1(_00371_),
    .C1(_00372_),
    .X(_01361_));
 sky130_fd_sc_hd__a211o_1 _08461_ (.A1(_00371_),
    .A2(_00372_),
    .B1(_00836_),
    .C1(_00837_),
    .X(_01362_));
 sky130_fd_sc_hd__o21a_1 _08462_ (.A1(_00832_),
    .A2(_01361_),
    .B1(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__a32o_1 _08463_ (.A1(net235),
    .A2(net249),
    .A3(_00828_),
    .B1(_00827_),
    .B2(_06383_),
    .X(_01364_));
 sky130_fd_sc_hd__clkbuf_4 _08464_ (.A(net206),
    .X(_01365_));
 sky130_fd_sc_hd__and4_1 _08465_ (.A(net235),
    .B(net208),
    .C(net250),
    .D(_01365_),
    .X(_01366_));
 sky130_fd_sc_hd__buf_2 _08466_ (.A(net250),
    .X(_01367_));
 sky130_fd_sc_hd__a22oi_1 _08467_ (.A1(net235),
    .A2(_01367_),
    .B1(_01365_),
    .B2(net208),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _08468_ (.A(_01366_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__and2_1 _08469_ (.A(_01364_),
    .B(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__nor2_1 _08470_ (.A(_01364_),
    .B(_01369_),
    .Y(_01371_));
 sky130_fd_sc_hd__or2_1 _08471_ (.A(_01370_),
    .B(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__xnor2_1 _08472_ (.A(_01363_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__xor2_1 _08473_ (.A(_00811_),
    .B(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__xnor2_1 _08474_ (.A(_00842_),
    .B(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__or2_1 _08475_ (.A(_01360_),
    .B(_01375_),
    .X(_01376_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(_01360_),
    .B(_01375_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _08477_ (.A(_01376_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__and2_1 _08478_ (.A(_00844_),
    .B(_00860_),
    .X(_01379_));
 sky130_fd_sc_hd__a22o_1 _08479_ (.A1(_06384_),
    .A2(_06383_),
    .B1(_00366_),
    .B2(_05980_),
    .X(_01380_));
 sky130_fd_sc_hd__nand4_4 _08480_ (.A(_05980_),
    .B(_06384_),
    .C(_06383_),
    .D(_00366_),
    .Y(_01381_));
 sky130_fd_sc_hd__a22o_1 _08481_ (.A1(_03853_),
    .A2(_00830_),
    .B1(_01380_),
    .B2(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__nand4_2 _08482_ (.A(_03853_),
    .B(_00830_),
    .C(_01380_),
    .D(_01381_),
    .Y(_01383_));
 sky130_fd_sc_hd__and2_1 _08483_ (.A(_01382_),
    .B(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_4 _08484_ (.A(net240),
    .X(_01385_));
 sky130_fd_sc_hd__and4_1 _08485_ (.A(_02492_),
    .B(_03864_),
    .C(_00834_),
    .D(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__a22o_1 _08486_ (.A1(_03864_),
    .A2(net240),
    .B1(net241),
    .B2(_02492_),
    .X(_01387_));
 sky130_fd_sc_hd__nand4_1 _08487_ (.A(_02492_),
    .B(_03864_),
    .C(net240),
    .D(net241),
    .Y(_01388_));
 sky130_fd_sc_hd__and2_1 _08488_ (.A(net246),
    .B(_00834_),
    .X(_01389_));
 sky130_fd_sc_hd__a21o_1 _08489_ (.A1(_01387_),
    .A2(_01388_),
    .B1(_01389_),
    .X(_01390_));
 sky130_fd_sc_hd__nand3_1 _08490_ (.A(_01387_),
    .B(_01388_),
    .C(_01389_),
    .Y(_01391_));
 sky130_fd_sc_hd__o211ai_1 _08491_ (.A1(_01386_),
    .A2(_00837_),
    .B1(_01390_),
    .C1(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__a211o_1 _08492_ (.A1(_01390_),
    .A2(_01391_),
    .B1(_01386_),
    .C1(_00837_),
    .X(_01393_));
 sky130_fd_sc_hd__nand2_1 _08493_ (.A(_01392_),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__xnor2_2 _08494_ (.A(_01384_),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__a21bo_1 _08495_ (.A1(_00845_),
    .A2(_00847_),
    .B1_N(_00846_),
    .X(_01396_));
 sky130_fd_sc_hd__clkbuf_4 _08496_ (.A(net13),
    .X(_01397_));
 sky130_fd_sc_hd__a22o_1 _08497_ (.A1(_03820_),
    .A2(_00821_),
    .B1(_01397_),
    .B2(net252),
    .X(_01398_));
 sky130_fd_sc_hd__nand4_1 _08498_ (.A(_03820_),
    .B(net252),
    .C(_00821_),
    .D(_01397_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(_01398_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__xnor2_2 _08500_ (.A(_01396_),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__xnor2_2 _08501_ (.A(_00824_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__xnor2_2 _08502_ (.A(_01395_),
    .B(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__inv_2 _08503_ (.A(_00852_),
    .Y(_01404_));
 sky130_fd_sc_hd__a21bo_1 _08504_ (.A1(_00355_),
    .A2(_01404_),
    .B1_N(_00854_),
    .X(_01405_));
 sky130_fd_sc_hd__a22o_1 _08505_ (.A1(net255),
    .A2(net9),
    .B1(net2),
    .B2(net8),
    .X(_01406_));
 sky130_fd_sc_hd__nand4_2 _08506_ (.A(_05882_),
    .B(_06375_),
    .C(_06368_),
    .D(net2),
    .Y(_01407_));
 sky130_fd_sc_hd__a22o_1 _08507_ (.A1(_05914_),
    .A2(_00822_),
    .B1(_01406_),
    .B2(_01407_),
    .X(_01408_));
 sky130_fd_sc_hd__nand4_1 _08508_ (.A(_05914_),
    .B(_00822_),
    .C(_01406_),
    .D(_01407_),
    .Y(_01409_));
 sky130_fd_sc_hd__clkbuf_4 _08509_ (.A(net4),
    .X(_01410_));
 sky130_fd_sc_hd__a22o_1 _08510_ (.A1(_03798_),
    .A2(_00850_),
    .B1(_01410_),
    .B2(_02470_),
    .X(_01411_));
 sky130_fd_sc_hd__and4_2 _08511_ (.A(net6),
    .B(_03798_),
    .C(net3),
    .D(net4),
    .X(_01412_));
 sky130_fd_sc_hd__xnor2_1 _08512_ (.A(_00852_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__and4_1 _08513_ (.A(_01408_),
    .B(_01409_),
    .C(_01411_),
    .D(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__a22oi_2 _08514_ (.A1(_01408_),
    .A2(_01409_),
    .B1(_01411_),
    .B2(_01413_),
    .Y(_01415_));
 sky130_fd_sc_hd__or3b_1 _08515_ (.A(_01414_),
    .B(_01415_),
    .C_N(_00876_),
    .X(_01416_));
 sky130_fd_sc_hd__o21bai_1 _08516_ (.A1(_01414_),
    .A2(_01415_),
    .B1_N(_00876_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand3_1 _08517_ (.A(_01405_),
    .B(_01416_),
    .C(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__a21o_1 _08518_ (.A1(_01416_),
    .A2(_01417_),
    .B1(_01405_),
    .X(_01419_));
 sky130_fd_sc_hd__a21o_1 _08519_ (.A1(_00857_),
    .A2(_00859_),
    .B1(_00856_),
    .X(_01420_));
 sky130_fd_sc_hd__and3_1 _08520_ (.A(_01418_),
    .B(_01419_),
    .C(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__a21oi_1 _08521_ (.A1(_01418_),
    .A2(_01419_),
    .B1(_01420_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _08522_ (.A(_01421_),
    .B(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__xor2_1 _08523_ (.A(_01403_),
    .B(_01423_),
    .X(_01424_));
 sky130_fd_sc_hd__o21a_1 _08524_ (.A1(_01379_),
    .A2(_00862_),
    .B1(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__nor3_1 _08525_ (.A(_01379_),
    .B(_00862_),
    .C(_01424_),
    .Y(_01426_));
 sky130_fd_sc_hd__or3_2 _08526_ (.A(_01378_),
    .B(_01425_),
    .C(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__o21ai_1 _08527_ (.A1(_01425_),
    .A2(_01426_),
    .B1(_01378_),
    .Y(_01428_));
 sky130_fd_sc_hd__and2_2 _08528_ (.A(_01427_),
    .B(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_00891_),
    .B(_00893_),
    .Y(_01430_));
 sky130_fd_sc_hd__a21bo_1 _08530_ (.A1(_00936_),
    .A2(_00948_),
    .B1_N(_00935_),
    .X(_01431_));
 sky130_fd_sc_hd__nand2_1 _08531_ (.A(_00887_),
    .B(_00889_),
    .Y(_01432_));
 sky130_fd_sc_hd__a21bo_1 _08532_ (.A1(_00880_),
    .A2(_00881_),
    .B1_N(_00882_),
    .X(_01433_));
 sky130_fd_sc_hd__clkbuf_4 _08533_ (.A(net65),
    .X(_01434_));
 sky130_fd_sc_hd__a22o_1 _08534_ (.A1(net52),
    .A2(_00397_),
    .B1(net64),
    .B2(net51),
    .X(_01435_));
 sky130_fd_sc_hd__nand4_2 _08535_ (.A(_03732_),
    .B(_05750_),
    .C(_00397_),
    .D(_00872_),
    .Y(_01436_));
 sky130_fd_sc_hd__a22o_1 _08536_ (.A1(_02580_),
    .A2(_01434_),
    .B1(_01435_),
    .B2(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__nand4_1 _08537_ (.A(_02580_),
    .B(_01434_),
    .C(_01435_),
    .D(_01436_),
    .Y(_01438_));
 sky130_fd_sc_hd__and3_1 _08538_ (.A(_01433_),
    .B(_01437_),
    .C(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__a21o_1 _08539_ (.A1(_01437_),
    .A2(_01438_),
    .B1(_01433_),
    .X(_01440_));
 sky130_fd_sc_hd__and2b_1 _08540_ (.A_N(_01439_),
    .B(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__xnor2_2 _08541_ (.A(_00874_),
    .B(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__buf_2 _08542_ (.A(net83),
    .X(_01443_));
 sky130_fd_sc_hd__buf_2 _08543_ (.A(net57),
    .X(_01444_));
 sky130_fd_sc_hd__a22oi_1 _08544_ (.A1(net68),
    .A2(_01443_),
    .B1(_01444_),
    .B2(net59),
    .Y(_01445_));
 sky130_fd_sc_hd__and4_1 _08545_ (.A(net68),
    .B(net59),
    .C(_01443_),
    .D(_01444_),
    .X(_01446_));
 sky130_fd_sc_hd__nor2_1 _08546_ (.A(_01445_),
    .B(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(_06343_),
    .B(_06347_),
    .Y(_01448_));
 sky130_fd_sc_hd__and3_1 _08548_ (.A(_03743_),
    .B(_05761_),
    .C(net54),
    .X(_01449_));
 sky130_fd_sc_hd__a22o_1 _08549_ (.A1(_05761_),
    .A2(net54),
    .B1(net55),
    .B2(_03743_),
    .X(_01450_));
 sky130_fd_sc_hd__a21bo_1 _08550_ (.A1(_00879_),
    .A2(_01449_),
    .B1_N(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__xor2_1 _08551_ (.A(_01448_),
    .B(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(_01447_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_1 _08553_ (.A(_00885_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__xor2_2 _08554_ (.A(_01442_),
    .B(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__and2_1 _08555_ (.A(_00425_),
    .B(_00946_),
    .X(_01456_));
 sky130_fd_sc_hd__xor2_2 _08556_ (.A(_01455_),
    .B(_01456_),
    .X(_01457_));
 sky130_fd_sc_hd__xnor2_2 _08557_ (.A(_01432_),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__xor2_2 _08558_ (.A(_01431_),
    .B(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__xnor2_2 _08559_ (.A(_01430_),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__and3_1 _08560_ (.A(_00869_),
    .B(_00893_),
    .C(_00894_),
    .X(_01461_));
 sky130_fd_sc_hd__a21oi_2 _08561_ (.A1(_00403_),
    .A2(_00896_),
    .B1(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__xnor2_2 _08562_ (.A(_01460_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__xor2_2 _08563_ (.A(_01429_),
    .B(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__xnor2_2 _08564_ (.A(_01358_),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__xnor2_2 _08565_ (.A(_01357_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__a31oi_2 _08566_ (.A1(net307),
    .A2(_00460_),
    .A3(_00965_),
    .B1(_00967_),
    .Y(_01467_));
 sky130_fd_sc_hd__and2_1 _08567_ (.A(_00526_),
    .B(_01017_),
    .X(_01468_));
 sky130_fd_sc_hd__or2_1 _08568_ (.A(_00939_),
    .B(_00942_),
    .X(_01469_));
 sky130_fd_sc_hd__a22oi_1 _08569_ (.A1(net71),
    .A2(_06410_),
    .B1(_00421_),
    .B2(_05498_),
    .Y(_01470_));
 sky130_fd_sc_hd__and4_1 _08570_ (.A(net70),
    .B(net71),
    .C(net80),
    .D(net81),
    .X(_01471_));
 sky130_fd_sc_hd__o2bb2a_1 _08571_ (.A1_N(_03579_),
    .A2_N(_00937_),
    .B1(_01470_),
    .B2(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__and4bb_1 _08572_ (.A_N(_01470_),
    .B_N(_01471_),
    .C(_03579_),
    .D(net82),
    .X(_01473_));
 sky130_fd_sc_hd__a211o_1 _08573_ (.A1(_00913_),
    .A2(_00915_),
    .B1(_01472_),
    .C1(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__o211ai_2 _08574_ (.A1(_01472_),
    .A2(_01473_),
    .B1(_00913_),
    .C1(_00915_),
    .Y(_01475_));
 sky130_fd_sc_hd__nand3_2 _08575_ (.A(_01469_),
    .B(_01474_),
    .C(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__a21o_1 _08576_ (.A1(_01474_),
    .A2(_01475_),
    .B1(_01469_),
    .X(_01477_));
 sky130_fd_sc_hd__and3_1 _08577_ (.A(_00917_),
    .B(_01476_),
    .C(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__a21oi_1 _08578_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_00917_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor3_1 _08579_ (.A(_00943_),
    .B(_00941_),
    .C(_00942_),
    .Y(_01480_));
 sky130_fd_sc_hd__o21ai_1 _08580_ (.A1(_00423_),
    .A2(_01480_),
    .B1(_00944_),
    .Y(_01481_));
 sky130_fd_sc_hd__or3_4 _08581_ (.A(_01478_),
    .B(_01479_),
    .C(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__o21ai_2 _08582_ (.A1(_01478_),
    .A2(_01479_),
    .B1(_01481_),
    .Y(_01483_));
 sky130_fd_sc_hd__clkbuf_4 _08583_ (.A(net119),
    .X(_01484_));
 sky130_fd_sc_hd__a22oi_2 _08584_ (.A1(_03524_),
    .A2(_00910_),
    .B1(_01484_),
    .B2(_02646_),
    .Y(_01485_));
 sky130_fd_sc_hd__and4_1 _08585_ (.A(_03524_),
    .B(net103),
    .C(_00910_),
    .D(_01484_),
    .X(_01486_));
 sky130_fd_sc_hd__clkbuf_4 _08586_ (.A(net73),
    .X(_01487_));
 sky130_fd_sc_hd__buf_2 _08587_ (.A(net74),
    .X(_01488_));
 sky130_fd_sc_hd__a22o_1 _08588_ (.A1(_03590_),
    .A2(_01487_),
    .B1(_01488_),
    .B2(_02657_),
    .X(_01489_));
 sky130_fd_sc_hd__nand4_2 _08589_ (.A(_02657_),
    .B(_03590_),
    .C(_01487_),
    .D(_01488_),
    .Y(_01490_));
 sky130_fd_sc_hd__a22o_1 _08590_ (.A1(_05520_),
    .A2(_00431_),
    .B1(_01489_),
    .B2(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__nand4_2 _08591_ (.A(_05520_),
    .B(_00431_),
    .C(_01489_),
    .D(_01490_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _08592_ (.A(_01491_),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor3_1 _08593_ (.A(_01485_),
    .B(_01486_),
    .C(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__o21a_1 _08594_ (.A1(_01485_),
    .A2(_01486_),
    .B1(_01493_),
    .X(_01495_));
 sky130_fd_sc_hd__nor2_1 _08595_ (.A(_01494_),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _08596_ (.A(_00922_),
    .B(_00924_),
    .Y(_01497_));
 sky130_fd_sc_hd__and4_1 _08597_ (.A(net113),
    .B(net114),
    .C(_00454_),
    .D(_00956_),
    .X(_01498_));
 sky130_fd_sc_hd__a22o_1 _08598_ (.A1(net106),
    .A2(net116),
    .B1(net107),
    .B2(net115),
    .X(_01499_));
 sky130_fd_sc_hd__nand4_2 _08599_ (.A(_05444_),
    .B(net106),
    .C(net116),
    .D(net107),
    .Y(_01500_));
 sky130_fd_sc_hd__a22o_1 _08600_ (.A1(_05389_),
    .A2(_00438_),
    .B1(_01499_),
    .B2(_01500_),
    .X(_01501_));
 sky130_fd_sc_hd__nand4_2 _08601_ (.A(_05389_),
    .B(_00438_),
    .C(_01499_),
    .D(_01500_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand3_1 _08602_ (.A(_01498_),
    .B(_01501_),
    .C(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__a21o_1 _08603_ (.A1(_01501_),
    .A2(_01502_),
    .B1(_01498_),
    .X(_01504_));
 sky130_fd_sc_hd__nand3_2 _08604_ (.A(_01497_),
    .B(_01503_),
    .C(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__a21o_1 _08605_ (.A1(_01503_),
    .A2(_01504_),
    .B1(_01497_),
    .X(_01506_));
 sky130_fd_sc_hd__a21bo_1 _08606_ (.A1(_00920_),
    .A2(_00926_),
    .B1_N(_00925_),
    .X(_01507_));
 sky130_fd_sc_hd__nand3_4 _08607_ (.A(_01505_),
    .B(_01506_),
    .C(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21o_1 _08608_ (.A1(_01505_),
    .A2(_01506_),
    .B1(_01507_),
    .X(_01509_));
 sky130_fd_sc_hd__nand3_4 _08609_ (.A(_01496_),
    .B(_01508_),
    .C(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21o_1 _08610_ (.A1(_01508_),
    .A2(_01509_),
    .B1(_01496_),
    .X(_01511_));
 sky130_fd_sc_hd__a21bo_1 _08611_ (.A1(_00919_),
    .A2(_00931_),
    .B1_N(_00930_),
    .X(_01512_));
 sky130_fd_sc_hd__nand3_4 _08612_ (.A(_01510_),
    .B(_01511_),
    .C(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__a21o_1 _08613_ (.A1(_01510_),
    .A2(_01511_),
    .B1(_01512_),
    .X(_01514_));
 sky130_fd_sc_hd__nand4_4 _08614_ (.A(_01482_),
    .B(_01483_),
    .C(_01513_),
    .D(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__a22o_1 _08615_ (.A1(_01482_),
    .A2(_01483_),
    .B1(_01513_),
    .B2(_01514_),
    .X(_01516_));
 sky130_fd_sc_hd__and3b_1 _08616_ (.A_N(_00959_),
    .B(_00960_),
    .C(_00476_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_1 _08617_ (.A(_00458_),
    .B(_00962_),
    .X(_01518_));
 sky130_fd_sc_hd__o21bai_2 _08618_ (.A1(_00984_),
    .A2(_00999_),
    .B1_N(_00998_),
    .Y(_01519_));
 sky130_fd_sc_hd__clkbuf_4 _08619_ (.A(net109),
    .X(_01520_));
 sky130_fd_sc_hd__a22oi_1 _08620_ (.A1(_03546_),
    .A2(_00956_),
    .B1(_01520_),
    .B2(_02635_),
    .Y(_01521_));
 sky130_fd_sc_hd__and4_1 _08621_ (.A(net113),
    .B(net114),
    .C(net108),
    .D(net109),
    .X(_01522_));
 sky130_fd_sc_hd__nor2_1 _08622_ (.A(_01521_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__clkbuf_4 _08623_ (.A(net180),
    .X(_01524_));
 sky130_fd_sc_hd__a22o_1 _08624_ (.A1(net100),
    .A2(net177),
    .B1(net178),
    .B2(net89),
    .X(_01525_));
 sky130_fd_sc_hd__nand4_1 _08625_ (.A(net89),
    .B(net100),
    .C(net177),
    .D(net178),
    .Y(_01526_));
 sky130_fd_sc_hd__a22oi_2 _08626_ (.A1(_02745_),
    .A2(_01524_),
    .B1(_01525_),
    .B2(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__and4_2 _08627_ (.A(net78),
    .B(net180),
    .C(_01525_),
    .D(_01526_),
    .X(_01528_));
 sky130_fd_sc_hd__or3_1 _08628_ (.A(_00955_),
    .B(_01527_),
    .C(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__o21ai_1 _08629_ (.A1(_01527_),
    .A2(_01528_),
    .B1(_00955_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand3_1 _08630_ (.A(_01523_),
    .B(_01529_),
    .C(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__a21o_1 _08631_ (.A1(_01529_),
    .A2(_01530_),
    .B1(_01523_),
    .X(_01532_));
 sky130_fd_sc_hd__nand3_1 _08632_ (.A(_00982_),
    .B(_01531_),
    .C(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__a21o_1 _08633_ (.A1(_01531_),
    .A2(_01532_),
    .B1(_00982_),
    .X(_01534_));
 sky130_fd_sc_hd__a21o_1 _08634_ (.A1(_01533_),
    .A2(_01534_),
    .B1(_00959_),
    .X(_01535_));
 sky130_fd_sc_hd__nand3_2 _08635_ (.A(_00959_),
    .B(_01533_),
    .C(_01534_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand3_4 _08636_ (.A(_01519_),
    .B(_01535_),
    .C(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__a21o_1 _08637_ (.A1(_01535_),
    .A2(_01536_),
    .B1(_01519_),
    .X(_01538_));
 sky130_fd_sc_hd__o211ai_4 _08638_ (.A1(_01517_),
    .A2(_01518_),
    .B1(_01537_),
    .C1(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__a211o_1 _08639_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01517_),
    .C1(_01518_),
    .X(_01540_));
 sky130_fd_sc_hd__or2b_1 _08640_ (.A(_00963_),
    .B_N(_00952_),
    .X(_01541_));
 sky130_fd_sc_hd__o21ai_1 _08641_ (.A1(_00463_),
    .A2(_00964_),
    .B1(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand3_2 _08642_ (.A(_01539_),
    .B(_01540_),
    .C(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_1 _08643_ (.A1(_01539_),
    .A2(_01540_),
    .B1(_01542_),
    .X(_01544_));
 sky130_fd_sc_hd__nand4_2 _08644_ (.A(_01515_),
    .B(_01516_),
    .C(_01543_),
    .D(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__a22o_1 _08645_ (.A1(_01515_),
    .A2(_01516_),
    .B1(_01543_),
    .B2(_01544_),
    .X(_01546_));
 sky130_fd_sc_hd__o211a_1 _08646_ (.A1(_01468_),
    .A2(_01019_),
    .B1(_01545_),
    .C1(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__a211oi_2 _08647_ (.A1(_01545_),
    .A2(_01546_),
    .B1(_01468_),
    .C1(_01019_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor3_1 _08648_ (.A(_01467_),
    .B(_01547_),
    .C(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__o21a_1 _08649_ (.A1(_01547_),
    .A2(_01548_),
    .B1(_01467_),
    .X(_01550_));
 sky130_fd_sc_hd__or2_1 _08650_ (.A(_00540_),
    .B(_01044_),
    .X(_01551_));
 sky130_fd_sc_hd__o21a_1 _08651_ (.A1(_01022_),
    .A2(_01045_),
    .B1(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__and3_1 _08652_ (.A(_05191_),
    .B(_00062_),
    .C(_00979_),
    .X(_01553_));
 sky130_fd_sc_hd__a22oi_1 _08653_ (.A1(_05202_),
    .A2(_00479_),
    .B1(_00985_),
    .B2(_03392_),
    .Y(_01554_));
 sky130_fd_sc_hd__and4_1 _08654_ (.A(net174),
    .B(net175),
    .C(_00479_),
    .D(_00985_),
    .X(_01555_));
 sky130_fd_sc_hd__nor2_1 _08655_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand2_1 _08656_ (.A(_00059_),
    .B(_00062_),
    .Y(_01557_));
 sky130_fd_sc_hd__xnor2_1 _08657_ (.A(_01556_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__o21a_1 _08658_ (.A1(_00978_),
    .A2(_01553_),
    .B1(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__nor3_1 _08659_ (.A(_00978_),
    .B(_01553_),
    .C(_01558_),
    .Y(_01560_));
 sky130_fd_sc_hd__or2_1 _08660_ (.A(_01559_),
    .B(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__buf_2 _08661_ (.A(net197),
    .X(_01562_));
 sky130_fd_sc_hd__buf_2 _08662_ (.A(net145),
    .X(_01563_));
 sky130_fd_sc_hd__a22oi_1 _08663_ (.A1(_02723_),
    .A2(_01562_),
    .B1(_01563_),
    .B2(net167),
    .Y(_01564_));
 sky130_fd_sc_hd__and4_1 _08664_ (.A(net182),
    .B(net167),
    .C(net197),
    .D(_01563_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _08665_ (.A(_01564_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__buf_2 _08666_ (.A(net196),
    .X(_01567_));
 sky130_fd_sc_hd__a22o_1 _08667_ (.A1(_00047_),
    .A2(_00989_),
    .B1(_00480_),
    .B2(net184),
    .X(_01568_));
 sky130_fd_sc_hd__nand4_1 _08668_ (.A(net184),
    .B(_00047_),
    .C(_00058_),
    .D(_00480_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand4_1 _08669_ (.A(_03337_),
    .B(_01567_),
    .C(_01568_),
    .D(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(net183),
    .A2(_01567_),
    .B1(_01568_),
    .B2(_01569_),
    .X(_01571_));
 sky130_fd_sc_hd__a21bo_1 _08671_ (.A1(_00988_),
    .A2(_00990_),
    .B1_N(_00991_),
    .X(_01572_));
 sky130_fd_sc_hd__nand3_1 _08672_ (.A(_01570_),
    .B(_01571_),
    .C(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__a21o_1 _08673_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01572_),
    .X(_01574_));
 sky130_fd_sc_hd__nand3_1 _08674_ (.A(_01566_),
    .B(_01573_),
    .C(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__a21o_1 _08675_ (.A1(_01573_),
    .A2(_01574_),
    .B1(_01566_),
    .X(_01576_));
 sky130_fd_sc_hd__o21bai_1 _08676_ (.A1(_00986_),
    .A2(_00995_),
    .B1_N(_00994_),
    .Y(_01577_));
 sky130_fd_sc_hd__and3_1 _08677_ (.A(_01575_),
    .B(_01576_),
    .C(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__a21oi_1 _08678_ (.A1(_01575_),
    .A2(_01576_),
    .B1(_01577_),
    .Y(_01579_));
 sky130_fd_sc_hd__or2_1 _08679_ (.A(_01578_),
    .B(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__xnor2_2 _08680_ (.A(_01561_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__and2b_1 _08681_ (.A_N(_01007_),
    .B(_01008_),
    .X(_01582_));
 sky130_fd_sc_hd__a31o_1 _08682_ (.A1(_02866_),
    .A2(_01023_),
    .A3(_01031_),
    .B1(_01030_),
    .X(_01583_));
 sky130_fd_sc_hd__clkbuf_4 _08683_ (.A(net188),
    .X(_01584_));
 sky130_fd_sc_hd__and3_1 _08684_ (.A(net191),
    .B(net192),
    .C(_01002_),
    .X(_01585_));
 sky130_fd_sc_hd__a22o_1 _08685_ (.A1(net192),
    .A2(net187),
    .B1(net188),
    .B2(net191),
    .X(_01586_));
 sky130_fd_sc_hd__a21bo_1 _08686_ (.A1(_01584_),
    .A2(_01585_),
    .B1_N(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__nand2_1 _08687_ (.A(net193),
    .B(_00489_),
    .Y(_01588_));
 sky130_fd_sc_hd__xnor2_1 _08688_ (.A(_01587_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__or2_1 _08689_ (.A(_01004_),
    .B(_01006_),
    .X(_01590_));
 sky130_fd_sc_hd__xor2_1 _08690_ (.A(_01589_),
    .B(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08691_ (.A(_01583_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__xnor2_1 _08692_ (.A(_01582_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__o21ai_1 _08693_ (.A1(_01013_),
    .A2(_01010_),
    .B1(_01011_),
    .Y(_01594_));
 sky130_fd_sc_hd__xnor2_1 _08694_ (.A(_01593_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__xor2_1 _08695_ (.A(_01581_),
    .B(_01595_),
    .X(_01596_));
 sky130_fd_sc_hd__xor2_1 _08696_ (.A(_01552_),
    .B(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__a22o_1 _08697_ (.A1(_01012_),
    .A2(_01014_),
    .B1(_01016_),
    .B2(_01001_),
    .X(_01598_));
 sky130_fd_sc_hd__or2b_1 _08698_ (.A(_01597_),
    .B_N(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__or2b_1 _08699_ (.A(_01598_),
    .B_N(_01597_),
    .X(_01600_));
 sky130_fd_sc_hd__nand2_1 _08700_ (.A(_01599_),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__and2_1 _08701_ (.A(_01033_),
    .B(_01043_),
    .X(_01602_));
 sky130_fd_sc_hd__buf_2 _08702_ (.A(net232),
    .X(_01603_));
 sky130_fd_sc_hd__a22oi_1 _08703_ (.A1(_03227_),
    .A2(_01023_),
    .B1(_01603_),
    .B2(net217),
    .Y(_01604_));
 sky130_fd_sc_hd__and4_1 _08704_ (.A(_03227_),
    .B(net217),
    .C(_01023_),
    .D(_01603_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _08705_ (.A(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__and4_1 _08706_ (.A(_04752_),
    .B(_04741_),
    .C(_00080_),
    .D(_00086_),
    .X(_01607_));
 sky130_fd_sc_hd__and4_1 _08707_ (.A(_03227_),
    .B(_00516_),
    .C(_01025_),
    .D(_01026_),
    .X(_01608_));
 sky130_fd_sc_hd__a22o_1 _08708_ (.A1(net220),
    .A2(net229),
    .B1(net221),
    .B2(net228),
    .X(_01609_));
 sky130_fd_sc_hd__nand4_4 _08709_ (.A(net228),
    .B(net220),
    .C(_00086_),
    .D(net221),
    .Y(_01610_));
 sky130_fd_sc_hd__nand4_2 _08710_ (.A(_04752_),
    .B(_00516_),
    .C(_01609_),
    .D(_01610_),
    .Y(_01611_));
 sky130_fd_sc_hd__a22o_1 _08711_ (.A1(_04752_),
    .A2(_00516_),
    .B1(_01609_),
    .B2(_01610_),
    .X(_01612_));
 sky130_fd_sc_hd__o211a_1 _08712_ (.A1(_01607_),
    .A2(_01608_),
    .B1(_01611_),
    .C1(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__a211o_1 _08713_ (.A1(_01611_),
    .A2(_01612_),
    .B1(_01607_),
    .C1(_01608_),
    .X(_01614_));
 sky130_fd_sc_hd__and2b_1 _08714_ (.A_N(_01613_),
    .B(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__xnor2_1 _08715_ (.A(_01606_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__clkbuf_4 _08716_ (.A(net224),
    .X(_01617_));
 sky130_fd_sc_hd__a22o_1 _08717_ (.A1(net227),
    .A2(_01034_),
    .B1(_01617_),
    .B2(net226),
    .X(_01618_));
 sky130_fd_sc_hd__nand4_2 _08718_ (.A(net226),
    .B(net227),
    .C(_01034_),
    .D(_01617_),
    .Y(_01619_));
 sky130_fd_sc_hd__and3_1 _08719_ (.A(_01053_),
    .B(_01618_),
    .C(_01619_),
    .X(_01620_));
 sky130_fd_sc_hd__a21o_1 _08720_ (.A1(_01618_),
    .A2(_01619_),
    .B1(_01053_),
    .X(_01621_));
 sky130_fd_sc_hd__and2b_1 _08721_ (.A_N(_01620_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_1 _08722_ (.A(_01037_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__xnor2_1 _08723_ (.A(_01616_),
    .B(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__xor2_1 _08724_ (.A(_01065_),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o21a_1 _08725_ (.A1(_01041_),
    .A2(_01602_),
    .B1(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__nor3_1 _08726_ (.A(_01041_),
    .B(_01602_),
    .C(_01625_),
    .Y(_01627_));
 sky130_fd_sc_hd__a21oi_1 _08727_ (.A1(_01054_),
    .A2(_01063_),
    .B1(_01061_),
    .Y(_01628_));
 sky130_fd_sc_hd__clkbuf_4 _08728_ (.A(net48),
    .X(_01629_));
 sky130_fd_sc_hd__nand2_1 _08729_ (.A(_02822_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__and3_1 _08730_ (.A(net33),
    .B(_04906_),
    .C(net47),
    .X(_01631_));
 sky130_fd_sc_hd__a22o_1 _08731_ (.A1(_04906_),
    .A2(net46),
    .B1(net47),
    .B2(net33),
    .X(_01632_));
 sky130_fd_sc_hd__a21bo_1 _08732_ (.A1(_00530_),
    .A2(_01631_),
    .B1_N(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__xor2_2 _08733_ (.A(_01630_),
    .B(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__a22o_1 _08734_ (.A1(net43),
    .A2(net37),
    .B1(net38),
    .B2(net42),
    .X(_01635_));
 sky130_fd_sc_hd__nand4_2 _08735_ (.A(_03194_),
    .B(_04862_),
    .C(_00543_),
    .D(_01068_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand4_1 _08736_ (.A(_00107_),
    .B(_00097_),
    .C(_01635_),
    .D(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__a22o_1 _08737_ (.A1(net36),
    .A2(_00097_),
    .B1(_01635_),
    .B2(_01636_),
    .X(_01638_));
 sky130_fd_sc_hd__a21bo_1 _08738_ (.A1(_01055_),
    .A2(_01056_),
    .B1_N(_01057_),
    .X(_01639_));
 sky130_fd_sc_hd__nand3_1 _08739_ (.A(_01637_),
    .B(_01638_),
    .C(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__a21o_1 _08740_ (.A1(_01637_),
    .A2(_01638_),
    .B1(_01639_),
    .X(_01641_));
 sky130_fd_sc_hd__and3_1 _08741_ (.A(_01634_),
    .B(_01640_),
    .C(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__a21oi_1 _08742_ (.A1(_01640_),
    .A2(_01641_),
    .B1(_01634_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor3b_1 _08743_ (.A(_01642_),
    .B(_01643_),
    .C_N(_01069_),
    .Y(_01644_));
 sky130_fd_sc_hd__o21ba_1 _08744_ (.A1(_01642_),
    .A2(_01643_),
    .B1_N(_01069_),
    .X(_01645_));
 sky130_fd_sc_hd__or3_2 _08745_ (.A(_01628_),
    .B(_01644_),
    .C(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__o21ai_1 _08746_ (.A1(_01644_),
    .A2(_01645_),
    .B1(_01628_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _08747_ (.A(_01646_),
    .B(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__inv_2 _08748_ (.A(_01089_),
    .Y(_01649_));
 sky130_fd_sc_hd__or3_4 _08749_ (.A(_01071_),
    .B(_01089_),
    .C(_01090_),
    .X(_01650_));
 sky130_fd_sc_hd__a31o_1 _08750_ (.A1(_02800_),
    .A2(_01072_),
    .A3(_01075_),
    .B1(_01074_),
    .X(_01651_));
 sky130_fd_sc_hd__buf_2 _08751_ (.A(net56),
    .X(_01652_));
 sky130_fd_sc_hd__clkbuf_4 _08752_ (.A(net39),
    .X(_01653_));
 sky130_fd_sc_hd__a22oi_1 _08753_ (.A1(_02800_),
    .A2(_01652_),
    .B1(_01653_),
    .B2(net41),
    .Y(_01654_));
 sky130_fd_sc_hd__and4_1 _08754_ (.A(_02800_),
    .B(net41),
    .C(_01652_),
    .D(_01653_),
    .X(_01655_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(_01654_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__and2_1 _08756_ (.A(_01651_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__nor2_1 _08757_ (.A(_01651_),
    .B(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _08758_ (.A(_01657_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(_03095_),
    .B(_01072_),
    .Y(_01660_));
 sky130_fd_sc_hd__and4_1 _08760_ (.A(net179),
    .B(_00549_),
    .C(_00109_),
    .D(_00544_),
    .X(_01661_));
 sky130_fd_sc_hd__a22o_1 _08761_ (.A1(_00549_),
    .A2(_00109_),
    .B1(_00544_),
    .B2(_04939_),
    .X(_01662_));
 sky130_fd_sc_hd__and2b_1 _08762_ (.A_N(_01661_),
    .B(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__xnor2_1 _08763_ (.A(_01660_),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__and2_1 _08764_ (.A(net12),
    .B(_00550_),
    .X(_01665_));
 sky130_fd_sc_hd__buf_2 _08765_ (.A(net212),
    .X(_01666_));
 sky130_fd_sc_hd__buf_2 _08766_ (.A(net223),
    .X(_01667_));
 sky130_fd_sc_hd__nand4_2 _08767_ (.A(_02789_),
    .B(_03106_),
    .C(_01666_),
    .D(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__a22o_1 _08768_ (.A1(_03106_),
    .A2(net212),
    .B1(net223),
    .B2(_02789_),
    .X(_01669_));
 sky130_fd_sc_hd__nand3_1 _08769_ (.A(_01665_),
    .B(_01668_),
    .C(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__a21o_1 _08770_ (.A1(_01668_),
    .A2(_01669_),
    .B1(_01665_),
    .X(_01671_));
 sky130_fd_sc_hd__a21bo_1 _08771_ (.A1(_01078_),
    .A2(_01080_),
    .B1_N(_01079_),
    .X(_01672_));
 sky130_fd_sc_hd__nand3_1 _08772_ (.A(_01670_),
    .B(_01671_),
    .C(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__a21o_1 _08773_ (.A1(_01670_),
    .A2(_01671_),
    .B1(_01672_),
    .X(_01674_));
 sky130_fd_sc_hd__nand3_1 _08774_ (.A(_01664_),
    .B(_01673_),
    .C(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__a21o_1 _08775_ (.A1(_01673_),
    .A2(_01674_),
    .B1(_01664_),
    .X(_01676_));
 sky130_fd_sc_hd__a21bo_1 _08776_ (.A1(_01077_),
    .A2(_01085_),
    .B1_N(_01084_),
    .X(_01677_));
 sky130_fd_sc_hd__nand3_2 _08777_ (.A(_01675_),
    .B(_01676_),
    .C(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__a21o_1 _08778_ (.A1(_01675_),
    .A2(_01676_),
    .B1(_01677_),
    .X(_01679_));
 sky130_fd_sc_hd__and3_2 _08779_ (.A(_01659_),
    .B(_01678_),
    .C(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__a21oi_2 _08780_ (.A1(_01678_),
    .A2(_01679_),
    .B1(_01659_),
    .Y(_01681_));
 sky130_fd_sc_hd__a211o_4 _08781_ (.A1(_01649_),
    .A2(_01650_),
    .B1(_01680_),
    .C1(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__o211ai_4 _08782_ (.A1(_01680_),
    .A2(_01681_),
    .B1(_01649_),
    .C1(_01650_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand3b_4 _08783_ (.A_N(_01648_),
    .B(_01682_),
    .C(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__a21bo_1 _08784_ (.A1(_01682_),
    .A2(_01683_),
    .B1_N(_01648_),
    .X(_01685_));
 sky130_fd_sc_hd__o211ai_4 _08785_ (.A1(_01093_),
    .A2(net300),
    .B1(_01684_),
    .C1(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__a211o_1 _08786_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01093_),
    .C1(net324),
    .X(_01687_));
 sky130_fd_sc_hd__or4bb_4 _08787_ (.A(_01626_),
    .B(_01627_),
    .C_N(_01686_),
    .D_N(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__a2bb2o_1 _08788_ (.A1_N(_01626_),
    .A2_N(_01627_),
    .B1(_01686_),
    .B2(_01687_),
    .X(_01689_));
 sky130_fd_sc_hd__o21bai_1 _08789_ (.A1(_01046_),
    .A2(_01098_),
    .B1_N(_01097_),
    .Y(_01690_));
 sky130_fd_sc_hd__and3_2 _08790_ (.A(_01688_),
    .B(_01689_),
    .C(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__a21oi_2 _08791_ (.A1(net310),
    .A2(_01689_),
    .B1(_01690_),
    .Y(_01692_));
 sky130_fd_sc_hd__or3_1 _08792_ (.A(_01601_),
    .B(_01691_),
    .C(_01692_),
    .X(_01693_));
 sky130_fd_sc_hd__o21ai_2 _08793_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01601_),
    .Y(_01694_));
 sky130_fd_sc_hd__o211a_1 _08794_ (.A1(_01101_),
    .A2(net294),
    .B1(_01693_),
    .C1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__a211o_1 _08795_ (.A1(_01693_),
    .A2(_01694_),
    .B1(_01101_),
    .C1(net323),
    .X(_01696_));
 sky130_fd_sc_hd__or4b_4 _08796_ (.A(_01549_),
    .B(_01550_),
    .C(_01695_),
    .D_N(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__o211ai_1 _08797_ (.A1(_01101_),
    .A2(net323),
    .B1(_01693_),
    .C1(_01694_),
    .Y(_01698_));
 sky130_fd_sc_hd__a2bb2o_1 _08798_ (.A1_N(_01549_),
    .A2_N(_01550_),
    .B1(_01698_),
    .B2(_01696_),
    .X(_01699_));
 sky130_fd_sc_hd__o211ai_4 _08799_ (.A1(_01105_),
    .A2(_01107_),
    .B1(_01697_),
    .C1(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__a211o_1 _08800_ (.A1(_01697_),
    .A2(_01699_),
    .B1(_01105_),
    .C1(net291),
    .X(_01701_));
 sky130_fd_sc_hd__nand3_2 _08801_ (.A(_01466_),
    .B(_01700_),
    .C(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(_01700_),
    .A2(_01701_),
    .B1(_01466_),
    .X(_01703_));
 sky130_fd_sc_hd__o211ai_4 _08803_ (.A1(_01109_),
    .A2(net290),
    .B1(_01702_),
    .C1(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__a211o_1 _08804_ (.A1(_01702_),
    .A2(_01703_),
    .B1(_01109_),
    .C1(net290),
    .X(_01705_));
 sky130_fd_sc_hd__nand4_2 _08805_ (.A(_01355_),
    .B(_01356_),
    .C(_01704_),
    .D(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__a22o_1 _08806_ (.A1(_01355_),
    .A2(_01356_),
    .B1(_01704_),
    .B2(_01705_),
    .X(_01707_));
 sky130_fd_sc_hd__o211ai_4 _08807_ (.A1(_01113_),
    .A2(net318),
    .B1(_01706_),
    .C1(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__a211o_1 _08808_ (.A1(_01706_),
    .A2(_01707_),
    .B1(_01113_),
    .C1(net318),
    .X(_01709_));
 sky130_fd_sc_hd__and3_2 _08809_ (.A(_01173_),
    .B(_01708_),
    .C(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__a21oi_2 _08810_ (.A1(_01708_),
    .A2(_01709_),
    .B1(_01173_),
    .Y(_01711_));
 sky130_fd_sc_hd__a211oi_4 _08811_ (.A1(_01117_),
    .A2(_01137_),
    .B1(_01710_),
    .C1(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__o211a_1 _08812_ (.A1(_01710_),
    .A2(_01711_),
    .B1(_01117_),
    .C1(_01137_),
    .X(_01713_));
 sky130_fd_sc_hd__nor3_1 _08813_ (.A(_01136_),
    .B(_01712_),
    .C(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__o21ai_1 _08814_ (.A1(_01712_),
    .A2(_01713_),
    .B1(_01136_),
    .Y(_01715_));
 sky130_fd_sc_hd__or2b_1 _08815_ (.A(_01714_),
    .B_N(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__o21bai_2 _08816_ (.A1(_00612_),
    .A2(_01122_),
    .B1_N(_01121_),
    .Y(_01717_));
 sky130_fd_sc_hd__xnor2_2 _08817_ (.A(_01716_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xnor2_1 _08818_ (.A(_01134_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__and2_1 _08819_ (.A(net282),
    .B(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__or2_1 _08820_ (.A(net282),
    .B(_01719_),
    .X(_01721_));
 sky130_fd_sc_hd__or2b_1 _08821_ (.A(_01720_),
    .B_N(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(net281),
    .B(_01128_),
    .Y(_01723_));
 sky130_fd_sc_hd__o21ai_1 _08823_ (.A1(_01129_),
    .A2(_01130_),
    .B1(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__xor2_1 _08824_ (.A(_01722_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__nor2_1 _08825_ (.A(_00166_),
    .B(_01725_),
    .Y(_00006_));
 sky130_fd_sc_hd__or2b_1 _08826_ (.A(_01138_),
    .B_N(_01172_),
    .X(_01726_));
 sky130_fd_sc_hd__o31ai_4 _08827_ (.A1(_01139_),
    .A2(_01169_),
    .A3(_01170_),
    .B1(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__inv_2 _08828_ (.A(_01708_),
    .Y(_01728_));
 sky130_fd_sc_hd__a21o_1 _08829_ (.A1(_01140_),
    .A2(_01167_),
    .B1(_01169_),
    .X(_01729_));
 sky130_fd_sc_hd__and2_1 _08830_ (.A(_01353_),
    .B(_01355_),
    .X(_01730_));
 sky130_fd_sc_hd__a41o_2 _08831_ (.A1(_06229_),
    .A2(_00177_),
    .A3(_00625_),
    .A4(_01166_),
    .B1(_01164_),
    .X(_01731_));
 sky130_fd_sc_hd__and2b_1 _08832_ (.A_N(_01279_),
    .B(_01280_),
    .X(_01732_));
 sky130_fd_sc_hd__o21ba_2 _08833_ (.A1(_01201_),
    .A2(_01281_),
    .B1_N(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__or2b_1 _08834_ (.A(_01200_),
    .B_N(_01176_),
    .X(_01734_));
 sky130_fd_sc_hd__a21bo_2 _08835_ (.A1(_01178_),
    .A2(_01199_),
    .B1_N(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__nor2_1 _08836_ (.A(_01189_),
    .B(_01191_),
    .Y(_01736_));
 sky130_fd_sc_hd__a22oi_2 _08837_ (.A1(_06227_),
    .A2(_00270_),
    .B1(_00171_),
    .B2(_06243_),
    .Y(_01737_));
 sky130_fd_sc_hd__and4_1 _08838_ (.A(_06243_),
    .B(_06227_),
    .C(_00270_),
    .D(_00171_),
    .X(_01738_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__nand2_1 _08840_ (.A(_06127_),
    .B(_00617_),
    .Y(_01740_));
 sky130_fd_sc_hd__xnor2_1 _08841_ (.A(_01739_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__xnor2_1 _08842_ (.A(_01736_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__or2_1 _08843_ (.A(_01145_),
    .B(_01148_),
    .X(_01743_));
 sky130_fd_sc_hd__xnor2_1 _08844_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__inv_2 _08845_ (.A(_01150_),
    .Y(_01745_));
 sky130_fd_sc_hd__o32a_1 _08846_ (.A1(_01143_),
    .A2(_01147_),
    .A3(_01148_),
    .B1(_01745_),
    .B2(_01151_),
    .X(_01746_));
 sky130_fd_sc_hd__xor2_1 _08847_ (.A(_01744_),
    .B(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__and2_1 _08848_ (.A(_04227_),
    .B(_01157_),
    .X(_01748_));
 sky130_fd_sc_hd__nor2_1 _08849_ (.A(_01747_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__and2_1 _08850_ (.A(_01747_),
    .B(_01748_),
    .X(_01750_));
 sky130_fd_sc_hd__or2_2 _08851_ (.A(_01749_),
    .B(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__o21ba_1 _08852_ (.A1(_01155_),
    .A2(_01158_),
    .B1_N(_01154_),
    .X(_01752_));
 sky130_fd_sc_hd__xor2_1 _08853_ (.A(_01751_),
    .B(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__buf_4 _08854_ (.A(net173),
    .X(_01754_));
 sky130_fd_sc_hd__and2_1 _08855_ (.A(_02328_),
    .B(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__or2_1 _08856_ (.A(_01753_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_2 _08857_ (.A(_01753_),
    .B(_01755_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_2 _08858_ (.A(_01756_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__xnor2_4 _08859_ (.A(_01735_),
    .B(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__xnor2_4 _08860_ (.A(_01161_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__xnor2_4 _08861_ (.A(_01733_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__xnor2_4 _08862_ (.A(_01731_),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__xnor2_2 _08863_ (.A(_01730_),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__xnor2_2 _08864_ (.A(_01729_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__inv_2 _08865_ (.A(_01704_),
    .Y(_01765_));
 sky130_fd_sc_hd__and4_1 _08866_ (.A(_01355_),
    .B(_01356_),
    .C(_01704_),
    .D(_01705_),
    .X(_01766_));
 sky130_fd_sc_hd__and2b_1 _08867_ (.A_N(_01349_),
    .B(_01351_),
    .X(_01767_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_01358_),
    .B(_01464_),
    .Y(_01768_));
 sky130_fd_sc_hd__or2b_1 _08869_ (.A(_01465_),
    .B_N(_01357_),
    .X(_01769_));
 sky130_fd_sc_hd__and2_1 _08870_ (.A(_01179_),
    .B(_01197_),
    .X(_01770_));
 sky130_fd_sc_hd__nor2_1 _08871_ (.A(_00651_),
    .B(_01198_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _08872_ (.A(_01240_),
    .B(_01241_),
    .Y(_01772_));
 sky130_fd_sc_hd__o21ba_1 _08873_ (.A1(_00648_),
    .A2(_01196_),
    .B1_N(_01194_),
    .X(_01773_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_00710_),
    .B(_01222_),
    .Y(_01774_));
 sky130_fd_sc_hd__and2_1 _08875_ (.A(_01185_),
    .B(_01192_),
    .X(_01775_));
 sky130_fd_sc_hd__o21ba_1 _08876_ (.A1(_00709_),
    .A2(_01206_),
    .B1_N(_01208_),
    .X(_01776_));
 sky130_fd_sc_hd__clkbuf_4 _08877_ (.A(net162),
    .X(_01777_));
 sky130_fd_sc_hd__a22o_1 _08878_ (.A1(net166),
    .A2(net163),
    .B1(net164),
    .B2(net165),
    .X(_01778_));
 sky130_fd_sc_hd__inv_2 _08879_ (.A(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__and4_1 _08880_ (.A(net165),
    .B(net166),
    .C(net163),
    .D(net164),
    .X(_01780_));
 sky130_fd_sc_hd__o2bb2a_1 _08881_ (.A1_N(_06130_),
    .A2_N(_01777_),
    .B1(_01779_),
    .B2(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__and4b_1 _08882_ (.A_N(_01780_),
    .B(_01777_),
    .C(net168),
    .D(_01778_),
    .X(_01782_));
 sky130_fd_sc_hd__nor2_1 _08883_ (.A(_01781_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__buf_2 _08884_ (.A(net31),
    .X(_01784_));
 sky130_fd_sc_hd__a22o_1 _08885_ (.A1(net17),
    .A2(net29),
    .B1(net30),
    .B2(net16),
    .X(_01785_));
 sky130_fd_sc_hd__inv_2 _08886_ (.A(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__and4_1 _08887_ (.A(net16),
    .B(_06138_),
    .C(_00647_),
    .D(_01181_),
    .X(_01787_));
 sky130_fd_sc_hd__o2bb2a_1 _08888_ (.A1_N(net15),
    .A2_N(_01784_),
    .B1(_01786_),
    .B2(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__and4b_1 _08889_ (.A_N(_01787_),
    .B(_01784_),
    .C(net15),
    .D(_01785_),
    .X(_01789_));
 sky130_fd_sc_hd__or2_2 _08890_ (.A(_01788_),
    .B(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__xnor2_2 _08891_ (.A(_01184_),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(_01783_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(_01776_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__xnor2_1 _08894_ (.A(_01775_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21o_1 _08895_ (.A1(_01774_),
    .A2(_01224_),
    .B1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__nand3_1 _08896_ (.A(_01774_),
    .B(_01224_),
    .C(_01794_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand3b_2 _08897_ (.A_N(_01773_),
    .B(_01795_),
    .C(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__a21bo_1 _08898_ (.A1(_01795_),
    .A2(_01796_),
    .B1_N(_01773_),
    .X(_01798_));
 sky130_fd_sc_hd__o211ai_4 _08899_ (.A1(_01772_),
    .A2(_01243_),
    .B1(_01797_),
    .C1(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__a211o_1 _08900_ (.A1(_01797_),
    .A2(_01798_),
    .B1(_01772_),
    .C1(_01243_),
    .X(_01800_));
 sky130_fd_sc_hd__o211ai_4 _08901_ (.A1(_01770_),
    .A2(_01771_),
    .B1(_01799_),
    .C1(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__a211o_1 _08902_ (.A1(_01799_),
    .A2(_01800_),
    .B1(_01770_),
    .C1(_01771_),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_1 _08903_ (.A(_01245_),
    .B(_01278_),
    .Y(_01803_));
 sky130_fd_sc_hd__and2_1 _08904_ (.A(_01227_),
    .B(_01239_),
    .X(_01804_));
 sky130_fd_sc_hd__or2b_1 _08905_ (.A(_01259_),
    .B_N(_01260_),
    .X(_01805_));
 sky130_fd_sc_hd__o31a_1 _08906_ (.A1(_01252_),
    .A2(_01253_),
    .A3(_01261_),
    .B1(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(_01231_),
    .B(_01233_),
    .Y(_01807_));
 sky130_fd_sc_hd__a22o_1 _08908_ (.A1(_06254_),
    .A2(net91),
    .B1(net92),
    .B2(_04413_),
    .X(_01808_));
 sky130_fd_sc_hd__nand4_1 _08909_ (.A(_04424_),
    .B(_06134_),
    .C(_00672_),
    .D(net92),
    .Y(_01809_));
 sky130_fd_sc_hd__a22oi_1 _08910_ (.A1(_06253_),
    .A2(_00200_),
    .B1(_01808_),
    .B2(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__and4_1 _08911_ (.A(_06253_),
    .B(_00200_),
    .C(_01808_),
    .D(_01809_),
    .X(_01811_));
 sky130_fd_sc_hd__nor2_1 _08912_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__xnor2_1 _08913_ (.A(_01253_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _08914_ (.A(_01807_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__xnor2_1 _08915_ (.A(_01806_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__xor2_1 _08916_ (.A(_01234_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__o21a_1 _08917_ (.A1(_01237_),
    .A2(_01804_),
    .B1(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__nor3_1 _08918_ (.A(_01237_),
    .B(_01804_),
    .C(_01816_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(_01203_),
    .B(_01205_),
    .Y(_01819_));
 sky130_fd_sc_hd__a22oi_1 _08920_ (.A1(net27),
    .A2(net19),
    .B1(net20),
    .B2(net26),
    .Y(_01820_));
 sky130_fd_sc_hd__and4_1 _08921_ (.A(net26),
    .B(net27),
    .C(net19),
    .D(net20),
    .X(_01821_));
 sky130_fd_sc_hd__o2bb2a_1 _08922_ (.A1_N(_06261_),
    .A2_N(net28),
    .B1(_01820_),
    .B2(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__and4bb_1 _08923_ (.A_N(_01820_),
    .B_N(_01821_),
    .C(_06261_),
    .D(net28),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_1 _08924_ (.A(_01822_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__xnor2_1 _08925_ (.A(_01220_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__xnor2_1 _08926_ (.A(_01819_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__or2_1 _08927_ (.A(_00705_),
    .B(_01215_),
    .X(_01827_));
 sky130_fd_sc_hd__or3_1 _08928_ (.A(_01216_),
    .B(_01219_),
    .C(_01220_),
    .X(_01828_));
 sky130_fd_sc_hd__and2_1 _08929_ (.A(net25),
    .B(net21),
    .X(_01829_));
 sky130_fd_sc_hd__nand4_1 _08930_ (.A(net85),
    .B(net24),
    .C(net102),
    .D(net22),
    .Y(_01830_));
 sky130_fd_sc_hd__a22o_1 _08931_ (.A1(net85),
    .A2(net102),
    .B1(net22),
    .B2(net24),
    .X(_01831_));
 sky130_fd_sc_hd__nand2_1 _08932_ (.A(_01830_),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__xnor2_1 _08933_ (.A(_01829_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _08934_ (.A(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__buf_2 _08935_ (.A(net101),
    .X(_01835_));
 sky130_fd_sc_hd__a22oi_1 _08936_ (.A1(net88),
    .A2(_00238_),
    .B1(_00703_),
    .B2(net87),
    .Y(_01836_));
 sky130_fd_sc_hd__and4_1 _08937_ (.A(net87),
    .B(net88),
    .C(net98),
    .D(net99),
    .X(_01837_));
 sky130_fd_sc_hd__o2bb2a_1 _08938_ (.A1_N(net86),
    .A2_N(_01835_),
    .B1(_01836_),
    .B2(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__and4bb_1 _08939_ (.A_N(_01836_),
    .B_N(_01837_),
    .C(net86),
    .D(net101),
    .X(_01839_));
 sky130_fd_sc_hd__nor2_1 _08940_ (.A(_01838_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__or2_1 _08941_ (.A(_01212_),
    .B(_01214_),
    .X(_01841_));
 sky130_fd_sc_hd__xnor2_1 _08942_ (.A(_01840_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__xnor2_1 _08943_ (.A(_01834_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_1 _08944_ (.A1(_01827_),
    .A2(_01828_),
    .B1(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__nand3_1 _08945_ (.A(_01827_),
    .B(_01828_),
    .C(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand3_1 _08946_ (.A(_01826_),
    .B(_01844_),
    .C(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__a21o_1 _08947_ (.A1(_01844_),
    .A2(_01845_),
    .B1(_01826_),
    .X(_01847_));
 sky130_fd_sc_hd__and2_1 _08948_ (.A(_01846_),
    .B(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__nor3b_1 _08949_ (.A(_01817_),
    .B(_01818_),
    .C_N(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__o21ba_1 _08950_ (.A1(_01817_),
    .A2(_01818_),
    .B1_N(_01848_),
    .X(_01850_));
 sky130_fd_sc_hd__or2_1 _08951_ (.A(_01249_),
    .B(_01273_),
    .X(_01851_));
 sky130_fd_sc_hd__or2b_1 _08952_ (.A(_01274_),
    .B_N(_01248_),
    .X(_01852_));
 sky130_fd_sc_hd__or2_1 _08953_ (.A(_01263_),
    .B(_01271_),
    .X(_01853_));
 sky130_fd_sc_hd__o21a_1 _08954_ (.A1(_01262_),
    .A2(_01272_),
    .B1(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__a22oi_1 _08955_ (.A1(_04303_),
    .A2(net137),
    .B1(net138),
    .B2(net121),
    .Y(_01855_));
 sky130_fd_sc_hd__and4_1 _08956_ (.A(_04303_),
    .B(net121),
    .C(net137),
    .D(net138),
    .X(_01856_));
 sky130_fd_sc_hd__nor2_1 _08957_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__clkbuf_4 _08958_ (.A(net93),
    .X(_01858_));
 sky130_fd_sc_hd__nand2_1 _08959_ (.A(net94),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xnor2_1 _08960_ (.A(_01857_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__a22o_1 _08961_ (.A1(net133),
    .A2(net126),
    .B1(net135),
    .B2(net125),
    .X(_01861_));
 sky130_fd_sc_hd__nand4_1 _08962_ (.A(net125),
    .B(net133),
    .C(net126),
    .D(net135),
    .Y(_01862_));
 sky130_fd_sc_hd__a22o_1 _08963_ (.A1(_06152_),
    .A2(_00665_),
    .B1(_01861_),
    .B2(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__nand4_1 _08964_ (.A(_06152_),
    .B(_00665_),
    .C(_01861_),
    .D(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21bo_1 _08965_ (.A1(_01255_),
    .A2(_01258_),
    .B1_N(_01256_),
    .X(_01865_));
 sky130_fd_sc_hd__nand3_1 _08966_ (.A(_01863_),
    .B(_01864_),
    .C(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__a21o_1 _08967_ (.A1(_01863_),
    .A2(_01864_),
    .B1(_01865_),
    .X(_01867_));
 sky130_fd_sc_hd__and3_1 _08968_ (.A(_01860_),
    .B(_01866_),
    .C(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__a21oi_1 _08969_ (.A1(_01866_),
    .A2(_01867_),
    .B1(_01860_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _08970_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__and2b_1 _08971_ (.A_N(_01270_),
    .B(_01269_),
    .X(_01871_));
 sky130_fd_sc_hd__clkbuf_4 _08972_ (.A(net129),
    .X(_01872_));
 sky130_fd_sc_hd__a22o_1 _08973_ (.A1(_04314_),
    .A2(_01264_),
    .B1(_01872_),
    .B2(net130),
    .X(_01873_));
 sky130_fd_sc_hd__nand4_2 _08974_ (.A(_02218_),
    .B(_04314_),
    .C(_01264_),
    .D(_01872_),
    .Y(_01874_));
 sky130_fd_sc_hd__a22o_1 _08975_ (.A1(_06151_),
    .A2(_00677_),
    .B1(_01873_),
    .B2(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__nand4_1 _08976_ (.A(_06151_),
    .B(_00677_),
    .C(_01873_),
    .D(_01874_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand3_1 _08977_ (.A(_01290_),
    .B(_01875_),
    .C(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__a21o_1 _08978_ (.A1(_01875_),
    .A2(_01876_),
    .B1(_01290_),
    .X(_01878_));
 sky130_fd_sc_hd__o2bb2ai_1 _08979_ (.A1_N(_01264_),
    .A2_N(_01265_),
    .B1(_01267_),
    .B2(_01268_),
    .Y(_01879_));
 sky130_fd_sc_hd__a21o_1 _08980_ (.A1(_01877_),
    .A2(_01878_),
    .B1(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__nand3_1 _08981_ (.A(_01877_),
    .B(_01878_),
    .C(_01879_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand3_1 _08982_ (.A(_01871_),
    .B(_01880_),
    .C(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21o_1 _08983_ (.A1(_01880_),
    .A2(_01881_),
    .B1(_01871_),
    .X(_01883_));
 sky130_fd_sc_hd__and3_1 _08984_ (.A(_01870_),
    .B(_01882_),
    .C(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__a21oi_2 _08985_ (.A1(_01882_),
    .A2(_01883_),
    .B1(_01870_),
    .Y(_01885_));
 sky130_fd_sc_hd__a211oi_4 _08986_ (.A1(_01303_),
    .A2(_01305_),
    .B1(_01884_),
    .C1(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__o211a_1 _08987_ (.A1(_01884_),
    .A2(_01885_),
    .B1(_01303_),
    .C1(_01305_),
    .X(_01887_));
 sky130_fd_sc_hd__nor3_2 _08988_ (.A(_01854_),
    .B(_01886_),
    .C(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__o21a_1 _08989_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01854_),
    .X(_01889_));
 sky130_fd_sc_hd__a211o_1 _08990_ (.A1(_01851_),
    .A2(_01852_),
    .B1(_01888_),
    .C1(_01889_),
    .X(_01890_));
 sky130_fd_sc_hd__o211ai_2 _08991_ (.A1(_01888_),
    .A2(_01889_),
    .B1(_01851_),
    .C1(_01852_),
    .Y(_01891_));
 sky130_fd_sc_hd__or4bb_4 _08992_ (.A(_01849_),
    .B(_01850_),
    .C_N(_01890_),
    .D_N(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__a2bb2o_1 _08993_ (.A1_N(_01849_),
    .A2_N(_01850_),
    .B1(_01890_),
    .B2(_01891_),
    .X(_01893_));
 sky130_fd_sc_hd__o211ai_4 _08994_ (.A1(_01276_),
    .A2(_01803_),
    .B1(_01892_),
    .C1(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a211o_1 _08995_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_01276_),
    .C1(_01803_),
    .X(_01895_));
 sky130_fd_sc_hd__nand4_4 _08996_ (.A(_01801_),
    .B(_01802_),
    .C(_01894_),
    .D(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__a22o_2 _08997_ (.A1(_01801_),
    .A2(_01802_),
    .B1(_01894_),
    .B2(_01895_),
    .X(_01897_));
 sky130_fd_sc_hd__nor3_2 _08998_ (.A(_01284_),
    .B(_01345_),
    .C(_01346_),
    .Y(_01898_));
 sky130_fd_sc_hd__and2b_1 _08999_ (.A_N(_01341_),
    .B(_01343_),
    .X(_01899_));
 sky130_fd_sc_hd__inv_2 _09000_ (.A(_01425_),
    .Y(_01900_));
 sky130_fd_sc_hd__nor2_1 _09001_ (.A(_01337_),
    .B(_01339_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(_00842_),
    .B(_01374_),
    .Y(_01902_));
 sky130_fd_sc_hd__o21bai_2 _09003_ (.A1(_01317_),
    .A2(_01320_),
    .B1_N(_01318_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand4_2 _09004_ (.A(net199),
    .B(net148),
    .C(net216),
    .D(net147),
    .Y(_01904_));
 sky130_fd_sc_hd__a22o_1 _09005_ (.A1(net199),
    .A2(net216),
    .B1(net147),
    .B2(net148),
    .X(_01905_));
 sky130_fd_sc_hd__a22o_1 _09006_ (.A1(net149),
    .A2(net146),
    .B1(_01904_),
    .B2(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__nand4_1 _09007_ (.A(net149),
    .B(_01309_),
    .C(_01904_),
    .D(_01905_),
    .Y(_01907_));
 sky130_fd_sc_hd__and3_1 _09008_ (.A(_01903_),
    .B(_01906_),
    .C(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__a21o_1 _09009_ (.A1(_01906_),
    .A2(_01907_),
    .B1(_01903_),
    .X(_01909_));
 sky130_fd_sc_hd__and2b_1 _09010_ (.A_N(_01908_),
    .B(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__xnor2_1 _09011_ (.A(_01311_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__a22o_1 _09012_ (.A1(_06361_),
    .A2(net213),
    .B1(net214),
    .B2(_06077_),
    .X(_01912_));
 sky130_fd_sc_hd__nand4_1 _09013_ (.A(_06086_),
    .B(_06361_),
    .C(net213),
    .D(_00757_),
    .Y(_01913_));
 sky130_fd_sc_hd__and2_1 _09014_ (.A(_03941_),
    .B(net215),
    .X(_01914_));
 sky130_fd_sc_hd__a21oi_1 _09015_ (.A1(_01912_),
    .A2(_01913_),
    .B1(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__and3_1 _09016_ (.A(_01912_),
    .B(_01913_),
    .C(_01914_),
    .X(_01916_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(_01915_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__and4_1 _09018_ (.A(_04106_),
    .B(_06173_),
    .C(_00343_),
    .D(_00810_),
    .X(_01918_));
 sky130_fd_sc_hd__and4_1 _09019_ (.A(_06362_),
    .B(_06304_),
    .C(_01324_),
    .D(_01325_),
    .X(_01919_));
 sky130_fd_sc_hd__a22o_1 _09020_ (.A1(_06172_),
    .A2(net205),
    .B1(net206),
    .B2(net209),
    .X(_01920_));
 sky130_fd_sc_hd__nand4_2 _09021_ (.A(_04106_),
    .B(_06173_),
    .C(net205),
    .D(net206),
    .Y(_01921_));
 sky130_fd_sc_hd__and2_1 _09022_ (.A(net211),
    .B(net204),
    .X(_01922_));
 sky130_fd_sc_hd__a21o_1 _09023_ (.A1(_01920_),
    .A2(_01921_),
    .B1(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__nand3_1 _09024_ (.A(_01920_),
    .B(_01921_),
    .C(_01922_),
    .Y(_01924_));
 sky130_fd_sc_hd__o211ai_2 _09025_ (.A1(_01918_),
    .A2(_01919_),
    .B1(_01923_),
    .C1(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__a211o_1 _09026_ (.A1(_01923_),
    .A2(_01924_),
    .B1(_01918_),
    .C1(_01919_),
    .X(_01926_));
 sky130_fd_sc_hd__nand3_1 _09027_ (.A(_01917_),
    .B(_01925_),
    .C(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__a21o_1 _09028_ (.A1(_01925_),
    .A2(_01926_),
    .B1(_01917_),
    .X(_01928_));
 sky130_fd_sc_hd__a21bo_1 _09029_ (.A1(_01321_),
    .A2(_01329_),
    .B1_N(_01328_),
    .X(_01929_));
 sky130_fd_sc_hd__and3_1 _09030_ (.A(_01927_),
    .B(_01928_),
    .C(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__a21oi_1 _09031_ (.A1(_01927_),
    .A2(_01928_),
    .B1(_01929_),
    .Y(_01931_));
 sky130_fd_sc_hd__or3_2 _09032_ (.A(_01911_),
    .B(_01930_),
    .C(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__o21ai_2 _09033_ (.A1(_01930_),
    .A2(_01931_),
    .B1(_01911_),
    .Y(_01933_));
 sky130_fd_sc_hd__o211a_1 _09034_ (.A1(_01333_),
    .A2(_01335_),
    .B1(_01932_),
    .C1(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__a211oi_2 _09035_ (.A1(_01932_),
    .A2(_01933_),
    .B1(_01333_),
    .C1(_01335_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(_01299_),
    .B(_01301_),
    .Y(_01936_));
 sky130_fd_sc_hd__a21o_1 _09037_ (.A1(_00775_),
    .A2(_01314_),
    .B1(_01313_),
    .X(_01937_));
 sky130_fd_sc_hd__a22oi_2 _09038_ (.A1(_06177_),
    .A2(net153),
    .B1(net154),
    .B2(net140),
    .Y(_01938_));
 sky130_fd_sc_hd__and4_1 _09039_ (.A(net140),
    .B(_06177_),
    .C(net153),
    .D(net154),
    .X(_01939_));
 sky130_fd_sc_hd__nor2_1 _09040_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__nand2_1 _09041_ (.A(net139),
    .B(net155),
    .Y(_01941_));
 sky130_fd_sc_hd__xnor2_1 _09042_ (.A(_01940_),
    .B(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__a22o_1 _09043_ (.A1(net151),
    .A2(net143),
    .B1(net144),
    .B2(net150),
    .X(_01943_));
 sky130_fd_sc_hd__nand4_2 _09044_ (.A(_06171_),
    .B(net151),
    .C(net143),
    .D(_00774_),
    .Y(_01944_));
 sky130_fd_sc_hd__a22oi_2 _09045_ (.A1(_06311_),
    .A2(_01293_),
    .B1(_01943_),
    .B2(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__and4_2 _09046_ (.A(_06311_),
    .B(_01293_),
    .C(_01943_),
    .D(_01944_),
    .X(_01946_));
 sky130_fd_sc_hd__a211o_1 _09047_ (.A1(_01296_),
    .A2(_01298_),
    .B1(_01945_),
    .C1(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__o211ai_2 _09048_ (.A1(_01945_),
    .A2(_01946_),
    .B1(_01296_),
    .C1(_01298_),
    .Y(_01948_));
 sky130_fd_sc_hd__nand3_1 _09049_ (.A(_01942_),
    .B(_01947_),
    .C(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__a21o_1 _09050_ (.A1(_01947_),
    .A2(_01948_),
    .B1(_01942_),
    .X(_01950_));
 sky130_fd_sc_hd__and3_1 _09051_ (.A(_01937_),
    .B(_01949_),
    .C(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__a21o_1 _09052_ (.A1(_01949_),
    .A2(_01950_),
    .B1(_01937_),
    .X(_01952_));
 sky130_fd_sc_hd__or2b_1 _09053_ (.A(_01951_),
    .B_N(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_2 _09054_ (.A(_01936_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor3b_2 _09055_ (.A(_01934_),
    .B(_01935_),
    .C_N(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__o21ba_1 _09056_ (.A1(_01934_),
    .A2(_01935_),
    .B1_N(_01954_),
    .X(_01956_));
 sky130_fd_sc_hd__a211oi_2 _09057_ (.A1(_01902_),
    .A2(_01376_),
    .B1(_01955_),
    .C1(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__o211a_1 _09058_ (.A1(_01955_),
    .A2(_01956_),
    .B1(_01902_),
    .C1(_01376_),
    .X(_01958_));
 sky130_fd_sc_hd__nor3_2 _09059_ (.A(_01901_),
    .B(_01957_),
    .C(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__o21a_1 _09060_ (.A1(_01957_),
    .A2(_01958_),
    .B1(_01901_),
    .X(_01960_));
 sky130_fd_sc_hd__a211oi_4 _09061_ (.A1(_01900_),
    .A2(_01427_),
    .B1(_01959_),
    .C1(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__o211a_1 _09062_ (.A1(_01959_),
    .A2(_01960_),
    .B1(_01900_),
    .C1(_01427_),
    .X(_01962_));
 sky130_fd_sc_hd__or3_4 _09063_ (.A(_01899_),
    .B(_01961_),
    .C(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__o21ai_4 _09064_ (.A1(_01961_),
    .A2(_01962_),
    .B1(_01899_),
    .Y(_01964_));
 sky130_fd_sc_hd__o211ai_4 _09065_ (.A1(_01345_),
    .A2(_01898_),
    .B1(_01963_),
    .C1(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__a211o_1 _09066_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01345_),
    .C1(_01898_),
    .X(_01966_));
 sky130_fd_sc_hd__and4_1 _09067_ (.A(_01896_),
    .B(_01897_),
    .C(_01965_),
    .D(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__a22oi_2 _09068_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_01965_),
    .B2(_01966_),
    .Y(_01968_));
 sky130_fd_sc_hd__a211o_1 _09069_ (.A1(_01768_),
    .A2(_01769_),
    .B1(_01967_),
    .C1(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__o211ai_1 _09070_ (.A1(_01967_),
    .A2(_01968_),
    .B1(_01768_),
    .C1(_01769_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand3b_1 _09071_ (.A_N(_01767_),
    .B(_01969_),
    .C(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__a21bo_1 _09072_ (.A1(_01969_),
    .A2(_01970_),
    .B1_N(_01767_),
    .X(_01972_));
 sky130_fd_sc_hd__and2_1 _09073_ (.A(_01971_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__inv_2 _09074_ (.A(_01700_),
    .Y(_01974_));
 sky130_fd_sc_hd__and3_1 _09075_ (.A(_01466_),
    .B(_01700_),
    .C(_01701_),
    .X(_01975_));
 sky130_fd_sc_hd__and2b_1 _09076_ (.A_N(_01462_),
    .B(_01460_),
    .X(_01976_));
 sky130_fd_sc_hd__a21oi_1 _09077_ (.A1(_01429_),
    .A2(_01463_),
    .B1(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__inv_2 _09078_ (.A(_01547_),
    .Y(_01978_));
 sky130_fd_sc_hd__or3_1 _09079_ (.A(_01467_),
    .B(_01547_),
    .C(_01548_),
    .X(_01979_));
 sky130_fd_sc_hd__or2_1 _09080_ (.A(_01363_),
    .B(_01372_),
    .X(_01980_));
 sky130_fd_sc_hd__o21a_1 _09081_ (.A1(_00811_),
    .A2(_01373_),
    .B1(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__inv_2 _09082_ (.A(_01402_),
    .Y(_01982_));
 sky130_fd_sc_hd__and2_1 _09083_ (.A(_00824_),
    .B(_01401_),
    .X(_01983_));
 sky130_fd_sc_hd__a21o_1 _09084_ (.A1(_01395_),
    .A2(_01982_),
    .B1(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__a21bo_1 _09085_ (.A1(_01384_),
    .A2(_01393_),
    .B1_N(_01392_),
    .X(_01985_));
 sky130_fd_sc_hd__clkbuf_4 _09086_ (.A(net207),
    .X(_01986_));
 sky130_fd_sc_hd__buf_2 _09087_ (.A(net251),
    .X(_01987_));
 sky130_fd_sc_hd__a22oi_1 _09088_ (.A1(_03853_),
    .A2(net250),
    .B1(_01987_),
    .B2(net235),
    .Y(_01988_));
 sky130_fd_sc_hd__and4_1 _09089_ (.A(net236),
    .B(net235),
    .C(net250),
    .D(net251),
    .X(_01989_));
 sky130_fd_sc_hd__o2bb2a_1 _09090_ (.A1_N(net208),
    .A2_N(_01986_),
    .B1(_01988_),
    .B2(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__and4bb_1 _09091_ (.A_N(_01988_),
    .B_N(_01989_),
    .C(net208),
    .D(_01986_),
    .X(_01991_));
 sky130_fd_sc_hd__a211o_1 _09092_ (.A1(_01381_),
    .A2(_01383_),
    .B1(_01990_),
    .C1(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__o211ai_2 _09093_ (.A1(_01990_),
    .A2(_01991_),
    .B1(_01381_),
    .C1(_01383_),
    .Y(_01993_));
 sky130_fd_sc_hd__a21o_1 _09094_ (.A1(_01992_),
    .A2(_01993_),
    .B1(_01366_),
    .X(_01994_));
 sky130_fd_sc_hd__nand3_1 _09095_ (.A(_01366_),
    .B(_01992_),
    .C(_01993_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand3_1 _09096_ (.A(_01985_),
    .B(_01994_),
    .C(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__a21o_1 _09097_ (.A1(_01994_),
    .A2(_01995_),
    .B1(_01985_),
    .X(_01997_));
 sky130_fd_sc_hd__a21o_1 _09098_ (.A1(_01996_),
    .A2(_01997_),
    .B1(_01370_),
    .X(_01998_));
 sky130_fd_sc_hd__nand3_1 _09099_ (.A(_01370_),
    .B(_01996_),
    .C(_01997_),
    .Y(_01999_));
 sky130_fd_sc_hd__and3_2 _09100_ (.A(_01984_),
    .B(_01998_),
    .C(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__a21oi_1 _09101_ (.A1(_01998_),
    .A2(_01999_),
    .B1(_01984_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _09102_ (.A(_02000_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__xor2_2 _09103_ (.A(_01981_),
    .B(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__and3_1 _09104_ (.A(net238),
    .B(net247),
    .C(_00366_),
    .X(_02004_));
 sky130_fd_sc_hd__a22o_1 _09105_ (.A1(net247),
    .A2(_00834_),
    .B1(_00366_),
    .B2(net238),
    .X(_02005_));
 sky130_fd_sc_hd__a21bo_1 _09106_ (.A1(_00834_),
    .A2(_02004_),
    .B1_N(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_2 _09107_ (.A(_05980_),
    .B(_00830_),
    .Y(_02007_));
 sky130_fd_sc_hd__xnor2_4 _09108_ (.A(_02006_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__a22o_1 _09109_ (.A1(net244),
    .A2(net241),
    .B1(net242),
    .B2(_02492_),
    .X(_02009_));
 sky130_fd_sc_hd__nand4_1 _09110_ (.A(_02492_),
    .B(_03864_),
    .C(net241),
    .D(net242),
    .Y(_02010_));
 sky130_fd_sc_hd__and2_1 _09111_ (.A(net246),
    .B(net240),
    .X(_02011_));
 sky130_fd_sc_hd__a21o_1 _09112_ (.A1(_02009_),
    .A2(_02010_),
    .B1(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__nand3_1 _09113_ (.A(_02009_),
    .B(_02010_),
    .C(_02011_),
    .Y(_02013_));
 sky130_fd_sc_hd__a21bo_1 _09114_ (.A1(_01387_),
    .A2(_01389_),
    .B1_N(_01388_),
    .X(_02014_));
 sky130_fd_sc_hd__and3_1 _09115_ (.A(_02012_),
    .B(_02013_),
    .C(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a21oi_1 _09116_ (.A1(_02012_),
    .A2(_02013_),
    .B1(_02014_),
    .Y(_02016_));
 sky130_fd_sc_hd__or2_2 _09117_ (.A(_02015_),
    .B(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__xor2_4 _09118_ (.A(_02008_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__clkbuf_4 _09119_ (.A(net14),
    .X(_02019_));
 sky130_fd_sc_hd__a22o_1 _09120_ (.A1(net254),
    .A2(net11),
    .B1(net13),
    .B2(_03820_),
    .X(_02020_));
 sky130_fd_sc_hd__nand4_2 _09121_ (.A(_03820_),
    .B(_05914_),
    .C(_00821_),
    .D(net13),
    .Y(_02021_));
 sky130_fd_sc_hd__a22o_1 _09122_ (.A1(net252),
    .A2(_02019_),
    .B1(_02020_),
    .B2(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__nand4_2 _09123_ (.A(_02481_),
    .B(_02019_),
    .C(_02020_),
    .D(_02021_),
    .Y(_02023_));
 sky130_fd_sc_hd__and4_1 _09124_ (.A(_05882_),
    .B(_06375_),
    .C(_06368_),
    .D(_00357_),
    .X(_02024_));
 sky130_fd_sc_hd__and4_1 _09125_ (.A(_05914_),
    .B(_00822_),
    .C(_01406_),
    .D(_01407_),
    .X(_02025_));
 sky130_fd_sc_hd__a211oi_1 _09126_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_02024_),
    .C1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__o211a_1 _09127_ (.A1(_02024_),
    .A2(_02025_),
    .B1(_02022_),
    .C1(_02023_),
    .X(_02027_));
 sky130_fd_sc_hd__nor2_1 _09128_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__and4_1 _09129_ (.A(_03820_),
    .B(_02481_),
    .C(_00821_),
    .D(_01397_),
    .X(_02029_));
 sky130_fd_sc_hd__and3_1 _09130_ (.A(_01396_),
    .B(_01398_),
    .C(_01399_),
    .X(_02030_));
 sky130_fd_sc_hd__nor2_1 _09131_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__xnor2_2 _09132_ (.A(_02028_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_4 _09133_ (.A(_02018_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__o21bai_4 _09134_ (.A1(_01404_),
    .A2(_01412_),
    .B1_N(_01414_),
    .Y(_02034_));
 sky130_fd_sc_hd__a21oi_2 _09135_ (.A1(_00874_),
    .A2(_01440_),
    .B1(_01439_),
    .Y(_02035_));
 sky130_fd_sc_hd__a22o_1 _09136_ (.A1(_06368_),
    .A2(net2),
    .B1(_00850_),
    .B2(_05882_),
    .X(_02036_));
 sky130_fd_sc_hd__nand4_1 _09137_ (.A(_05882_),
    .B(_06368_),
    .C(_00357_),
    .D(_00850_),
    .Y(_02037_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(_02036_),
    .B(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__and2_1 _09139_ (.A(_06375_),
    .B(net10),
    .X(_02039_));
 sky130_fd_sc_hd__xor2_2 _09140_ (.A(_02038_),
    .B(_02039_),
    .X(_02040_));
 sky130_fd_sc_hd__a22oi_1 _09141_ (.A1(net50),
    .A2(net66),
    .B1(net5),
    .B2(_02470_),
    .Y(_02041_));
 sky130_fd_sc_hd__and4_1 _09142_ (.A(net50),
    .B(net6),
    .C(net66),
    .D(net5),
    .X(_02042_));
 sky130_fd_sc_hd__or2_1 _09143_ (.A(_02041_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__and2_1 _09144_ (.A(_03798_),
    .B(net4),
    .X(_02044_));
 sky130_fd_sc_hd__a21bo_1 _09145_ (.A1(_02470_),
    .A2(_00850_),
    .B1_N(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__xnor2_2 _09146_ (.A(_02043_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__xnor2_2 _09147_ (.A(_02040_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__xor2_2 _09148_ (.A(_02035_),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__xor2_2 _09149_ (.A(_02034_),
    .B(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__and2_1 _09150_ (.A(_01416_),
    .B(_01418_),
    .X(_02050_));
 sky130_fd_sc_hd__xnor2_2 _09151_ (.A(_02049_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__xor2_2 _09152_ (.A(_02033_),
    .B(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__a21oi_2 _09153_ (.A1(_01403_),
    .A2(_01423_),
    .B1(_01421_),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_2 _09154_ (.A(_02052_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__xnor2_2 _09155_ (.A(_02003_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__and2b_1 _09156_ (.A_N(_01458_),
    .B(_01431_),
    .X(_02056_));
 sky130_fd_sc_hd__and2b_1 _09157_ (.A_N(_01459_),
    .B(_01430_),
    .X(_02057_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_01455_),
    .B(_01456_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21bo_1 _09159_ (.A1(_01432_),
    .A2(_01457_),
    .B1_N(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__or2_1 _09160_ (.A(_00885_),
    .B(_01453_),
    .X(_02060_));
 sky130_fd_sc_hd__or2_1 _09161_ (.A(_01442_),
    .B(_01454_),
    .X(_02061_));
 sky130_fd_sc_hd__nand3_1 _09162_ (.A(_00917_),
    .B(_01476_),
    .C(_01477_),
    .Y(_02062_));
 sky130_fd_sc_hd__and2_1 _09163_ (.A(_01447_),
    .B(_01452_),
    .X(_02063_));
 sky130_fd_sc_hd__buf_2 _09164_ (.A(net84),
    .X(_02064_));
 sky130_fd_sc_hd__a22o_1 _09165_ (.A1(net69),
    .A2(net83),
    .B1(_02064_),
    .B2(net68),
    .X(_02065_));
 sky130_fd_sc_hd__nand4_1 _09166_ (.A(net69),
    .B(net68),
    .C(_01443_),
    .D(_02064_),
    .Y(_02066_));
 sky130_fd_sc_hd__and2_1 _09167_ (.A(net59),
    .B(net58),
    .X(_02067_));
 sky130_fd_sc_hd__a21o_1 _09168_ (.A1(_02065_),
    .A2(_02066_),
    .B1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nand3_1 _09169_ (.A(_02065_),
    .B(_02066_),
    .C(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand3_1 _09170_ (.A(_01446_),
    .B(_02068_),
    .C(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21o_1 _09171_ (.A1(_02068_),
    .A2(_02069_),
    .B1(_01446_),
    .X(_02071_));
 sky130_fd_sc_hd__and3_1 _09172_ (.A(net60),
    .B(net61),
    .C(net55),
    .X(_02072_));
 sky130_fd_sc_hd__a22o_1 _09173_ (.A1(net61),
    .A2(net55),
    .B1(net57),
    .B2(net60),
    .X(_02073_));
 sky130_fd_sc_hd__a21bo_1 _09174_ (.A1(_01444_),
    .A2(_02072_),
    .B1_N(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(_06347_),
    .B(_00387_),
    .Y(_02075_));
 sky130_fd_sc_hd__xor2_2 _09176_ (.A(_02074_),
    .B(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__a21o_1 _09177_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__nand3_1 _09178_ (.A(_02070_),
    .B(_02071_),
    .C(_02076_),
    .Y(_02078_));
 sky130_fd_sc_hd__and3_1 _09179_ (.A(_02063_),
    .B(_02077_),
    .C(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__a21oi_1 _09180_ (.A1(_02077_),
    .A2(_02078_),
    .B1(_02063_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _09181_ (.A(_01436_),
    .B(_01438_),
    .Y(_02081_));
 sky130_fd_sc_hd__a32o_1 _09182_ (.A1(_06343_),
    .A2(_06347_),
    .A3(_01450_),
    .B1(_01449_),
    .B2(_00879_),
    .X(_02082_));
 sky130_fd_sc_hd__a22o_1 _09183_ (.A1(net53),
    .A2(net63),
    .B1(net64),
    .B2(net52),
    .X(_02083_));
 sky130_fd_sc_hd__nand4_2 _09184_ (.A(_05750_),
    .B(net53),
    .C(_00397_),
    .D(_00872_),
    .Y(_02084_));
 sky130_fd_sc_hd__a22o_1 _09185_ (.A1(_03732_),
    .A2(_01434_),
    .B1(_02083_),
    .B2(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand4_1 _09186_ (.A(_03732_),
    .B(_01434_),
    .C(_02083_),
    .D(_02084_),
    .Y(_02086_));
 sky130_fd_sc_hd__and3_1 _09187_ (.A(_02082_),
    .B(_02085_),
    .C(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__a21o_1 _09188_ (.A1(_02085_),
    .A2(_02086_),
    .B1(_02082_),
    .X(_02088_));
 sky130_fd_sc_hd__or2b_1 _09189_ (.A(_02087_),
    .B_N(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__xnor2_1 _09190_ (.A(_02081_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor3b_1 _09191_ (.A(_02079_),
    .B(_02080_),
    .C_N(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__o21ba_1 _09192_ (.A1(_02079_),
    .A2(_02080_),
    .B1_N(_02090_),
    .X(_02092_));
 sky130_fd_sc_hd__a211oi_2 _09193_ (.A1(_02062_),
    .A2(_01482_),
    .B1(net305),
    .C1(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__o211a_1 _09194_ (.A1(net305),
    .A2(_02092_),
    .B1(_02062_),
    .C1(_01482_),
    .X(_02094_));
 sky130_fd_sc_hd__a211oi_2 _09195_ (.A1(_02060_),
    .A2(_02061_),
    .B1(_02093_),
    .C1(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__o211a_1 _09196_ (.A1(_02093_),
    .A2(_02094_),
    .B1(_02060_),
    .C1(_02061_),
    .X(_02096_));
 sky130_fd_sc_hd__a211o_1 _09197_ (.A1(_01513_),
    .A2(_01515_),
    .B1(_02095_),
    .C1(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__o211ai_2 _09198_ (.A1(_02095_),
    .A2(_02096_),
    .B1(_01513_),
    .C1(_01515_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand3_1 _09199_ (.A(_02059_),
    .B(_02097_),
    .C(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__a21o_1 _09200_ (.A1(_02097_),
    .A2(_02098_),
    .B1(_02059_),
    .X(_02100_));
 sky130_fd_sc_hd__o211ai_2 _09201_ (.A1(_02056_),
    .A2(_02057_),
    .B1(_02099_),
    .C1(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__a211o_1 _09202_ (.A1(_02099_),
    .A2(_02100_),
    .B1(_02056_),
    .C1(_02057_),
    .X(_02102_));
 sky130_fd_sc_hd__and3_1 _09203_ (.A(_02055_),
    .B(_02101_),
    .C(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__a21oi_1 _09204_ (.A1(_02101_),
    .A2(_02102_),
    .B1(_02055_),
    .Y(_02104_));
 sky130_fd_sc_hd__a211oi_2 _09205_ (.A1(_01978_),
    .A2(_01979_),
    .B1(_02103_),
    .C1(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__o211a_1 _09206_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_01978_),
    .C1(_01979_),
    .X(_02106_));
 sky130_fd_sc_hd__nor3_1 _09207_ (.A(_01977_),
    .B(_02105_),
    .C(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__o21a_1 _09208_ (.A1(_02105_),
    .A2(_02106_),
    .B1(_01977_),
    .X(_02108_));
 sky130_fd_sc_hd__nor2_2 _09209_ (.A(_02107_),
    .B(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__and4bb_1 _09210_ (.A_N(_01549_),
    .B_N(_01550_),
    .C(_01698_),
    .D(_01696_),
    .X(_02110_));
 sky130_fd_sc_hd__nand2_1 _09211_ (.A(_01543_),
    .B(_01545_),
    .Y(_02111_));
 sky130_fd_sc_hd__or2b_1 _09212_ (.A(_01552_),
    .B_N(_01596_),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(_01474_),
    .B(_01476_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _09214_ (.A(_01471_),
    .B(_01473_),
    .Y(_02114_));
 sky130_fd_sc_hd__a22o_1 _09215_ (.A1(net80),
    .A2(net72),
    .B1(net81),
    .B2(net71),
    .X(_02115_));
 sky130_fd_sc_hd__nand4_1 _09216_ (.A(_06424_),
    .B(_06410_),
    .C(net72),
    .D(_00421_),
    .Y(_02116_));
 sky130_fd_sc_hd__a22oi_2 _09217_ (.A1(_05498_),
    .A2(_00937_),
    .B1(_02115_),
    .B2(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__and4_1 _09218_ (.A(_05498_),
    .B(_00937_),
    .C(_02115_),
    .D(_02116_),
    .X(_02118_));
 sky130_fd_sc_hd__a211o_1 _09219_ (.A1(_01490_),
    .A2(_01492_),
    .B1(_02117_),
    .C1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__o211ai_1 _09220_ (.A1(_02117_),
    .A2(_02118_),
    .B1(_01490_),
    .C1(_01492_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand3b_1 _09221_ (.A_N(_02114_),
    .B(_02119_),
    .C(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__a21bo_1 _09222_ (.A1(_02119_),
    .A2(_02120_),
    .B1_N(_02114_),
    .X(_02122_));
 sky130_fd_sc_hd__and3_1 _09223_ (.A(_01494_),
    .B(_02121_),
    .C(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__a21o_1 _09224_ (.A1(_02121_),
    .A2(_02122_),
    .B1(_01494_),
    .X(_02124_));
 sky130_fd_sc_hd__or2b_1 _09225_ (.A(_02123_),
    .B_N(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__xnor2_2 _09226_ (.A(_02113_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__and3_1 _09227_ (.A(net76),
    .B(net77),
    .C(net74),
    .X(_02127_));
 sky130_fd_sc_hd__a22o_1 _09228_ (.A1(net77),
    .A2(net74),
    .B1(net75),
    .B2(net76),
    .X(_02128_));
 sky130_fd_sc_hd__a21bo_1 _09229_ (.A1(net75),
    .A2(_02127_),
    .B1_N(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_05520_),
    .B(_01487_),
    .Y(_02130_));
 sky130_fd_sc_hd__xor2_1 _09231_ (.A(_02129_),
    .B(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__clkbuf_4 _09232_ (.A(net120),
    .X(_02132_));
 sky130_fd_sc_hd__a22o_1 _09233_ (.A1(net105),
    .A2(net118),
    .B1(net119),
    .B2(net104),
    .X(_02133_));
 sky130_fd_sc_hd__nand4_2 _09234_ (.A(net104),
    .B(net105),
    .C(net118),
    .D(net119),
    .Y(_02134_));
 sky130_fd_sc_hd__a22o_1 _09235_ (.A1(net103),
    .A2(_02132_),
    .B1(_02133_),
    .B2(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__nand4_1 _09236_ (.A(net103),
    .B(_02132_),
    .C(_02133_),
    .D(_02134_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand3_1 _09237_ (.A(_01486_),
    .B(_02135_),
    .C(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__a21o_1 _09238_ (.A1(_02135_),
    .A2(_02136_),
    .B1(_01486_),
    .X(_02138_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(_02137_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__xnor2_1 _09240_ (.A(_02131_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _09241_ (.A(_01500_),
    .B(_01502_),
    .Y(_02141_));
 sky130_fd_sc_hd__a22o_1 _09242_ (.A1(net116),
    .A2(net107),
    .B1(net108),
    .B2(net115),
    .X(_02142_));
 sky130_fd_sc_hd__nand4_2 _09243_ (.A(net115),
    .B(net116),
    .C(net107),
    .D(net108),
    .Y(_02143_));
 sky130_fd_sc_hd__a22o_1 _09244_ (.A1(_06437_),
    .A2(net117),
    .B1(_02142_),
    .B2(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__nand4_2 _09245_ (.A(_06437_),
    .B(net117),
    .C(_02142_),
    .D(_02143_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand3_1 _09246_ (.A(_01522_),
    .B(_02144_),
    .C(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__a21o_1 _09247_ (.A1(_02144_),
    .A2(_02145_),
    .B1(_01522_),
    .X(_02147_));
 sky130_fd_sc_hd__nand3_1 _09248_ (.A(_02141_),
    .B(_02146_),
    .C(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__a21o_1 _09249_ (.A1(_02146_),
    .A2(_02147_),
    .B1(_02141_),
    .X(_02149_));
 sky130_fd_sc_hd__a21bo_1 _09250_ (.A1(_01497_),
    .A2(_01504_),
    .B1_N(_01503_),
    .X(_02150_));
 sky130_fd_sc_hd__nand3_1 _09251_ (.A(_02148_),
    .B(_02149_),
    .C(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__a21o_1 _09252_ (.A1(_02148_),
    .A2(_02149_),
    .B1(_02150_),
    .X(_02152_));
 sky130_fd_sc_hd__and3_2 _09253_ (.A(_02140_),
    .B(_02151_),
    .C(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__a21oi_2 _09254_ (.A1(_02151_),
    .A2(_02152_),
    .B1(_02140_),
    .Y(_02154_));
 sky130_fd_sc_hd__a211o_1 _09255_ (.A1(_01508_),
    .A2(_01510_),
    .B1(_02153_),
    .C1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__o211ai_4 _09256_ (.A1(_02153_),
    .A2(_02154_),
    .B1(_01508_),
    .C1(_01510_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand3_2 _09257_ (.A(_02126_),
    .B(_02155_),
    .C(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__a21o_1 _09258_ (.A1(_02155_),
    .A2(_02156_),
    .B1(_02126_),
    .X(_02158_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_01533_),
    .B(_01536_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand3_1 _09260_ (.A(_01575_),
    .B(_01576_),
    .C(_01577_),
    .Y(_02160_));
 sky130_fd_sc_hd__or3_1 _09261_ (.A(_01561_),
    .B(_01578_),
    .C(_01579_),
    .X(_02161_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(_01529_),
    .B(_01531_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(_03546_),
    .B(net109),
    .Y(_02163_));
 sky130_fd_sc_hd__clkbuf_4 _09264_ (.A(net110),
    .X(_02164_));
 sky130_fd_sc_hd__and3_1 _09265_ (.A(net78),
    .B(net113),
    .C(net181),
    .X(_02165_));
 sky130_fd_sc_hd__a22o_1 _09266_ (.A1(net78),
    .A2(net181),
    .B1(net110),
    .B2(net113),
    .X(_02166_));
 sky130_fd_sc_hd__a21bo_1 _09267_ (.A1(_02164_),
    .A2(_02165_),
    .B1_N(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__xor2_2 _09268_ (.A(_02163_),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__and4_1 _09269_ (.A(net89),
    .B(net100),
    .C(_00453_),
    .D(_00953_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _09270_ (.A1(net111),
    .A2(net177),
    .B1(net178),
    .B2(net100),
    .X(_02170_));
 sky130_fd_sc_hd__nand4_2 _09271_ (.A(net100),
    .B(net111),
    .C(_00453_),
    .D(_00953_),
    .Y(_02171_));
 sky130_fd_sc_hd__a22o_1 _09272_ (.A1(net89),
    .A2(_01524_),
    .B1(_02170_),
    .B2(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__nand4_2 _09273_ (.A(_03381_),
    .B(_01524_),
    .C(_02170_),
    .D(_02171_),
    .Y(_02173_));
 sky130_fd_sc_hd__o211ai_2 _09274_ (.A1(_02169_),
    .A2(_01528_),
    .B1(_02172_),
    .C1(_02173_),
    .Y(_02175_));
 sky130_fd_sc_hd__a211o_1 _09275_ (.A1(_02172_),
    .A2(_02173_),
    .B1(_02169_),
    .C1(_01528_),
    .X(_02176_));
 sky130_fd_sc_hd__nand3_2 _09276_ (.A(_02168_),
    .B(_02175_),
    .C(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__a21o_1 _09277_ (.A1(_02175_),
    .A2(_02176_),
    .B1(_02168_),
    .X(_02178_));
 sky130_fd_sc_hd__nand3_1 _09278_ (.A(_01559_),
    .B(_02177_),
    .C(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__a21o_1 _09279_ (.A1(_02177_),
    .A2(_02178_),
    .B1(_01559_),
    .X(_02180_));
 sky130_fd_sc_hd__and3_1 _09280_ (.A(_02162_),
    .B(_02179_),
    .C(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__a21oi_1 _09281_ (.A1(_02179_),
    .A2(_02180_),
    .B1(_02162_),
    .Y(_02182_));
 sky130_fd_sc_hd__a211o_1 _09282_ (.A1(_02160_),
    .A2(_02161_),
    .B1(_02181_),
    .C1(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__o211ai_2 _09283_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02160_),
    .C1(_02161_),
    .Y(_02184_));
 sky130_fd_sc_hd__and3_1 _09284_ (.A(_02159_),
    .B(_02183_),
    .C(_02184_),
    .X(_02186_));
 sky130_fd_sc_hd__a21oi_1 _09285_ (.A1(_02183_),
    .A2(_02184_),
    .B1(_02159_),
    .Y(_02187_));
 sky130_fd_sc_hd__a211o_1 _09286_ (.A1(_01537_),
    .A2(_01539_),
    .B1(_02186_),
    .C1(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__o211ai_2 _09287_ (.A1(_02186_),
    .A2(_02187_),
    .B1(_01537_),
    .C1(_01539_),
    .Y(_02189_));
 sky130_fd_sc_hd__and4_1 _09288_ (.A(_02157_),
    .B(_02158_),
    .C(_02188_),
    .D(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a22oi_2 _09289_ (.A1(_02157_),
    .A2(_02158_),
    .B1(_02188_),
    .B2(_02189_),
    .Y(_02191_));
 sky130_fd_sc_hd__a211o_1 _09290_ (.A1(_02112_),
    .A2(_01599_),
    .B1(_02190_),
    .C1(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__o211ai_2 _09291_ (.A1(_02190_),
    .A2(_02191_),
    .B1(_02112_),
    .C1(_01599_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand3_1 _09292_ (.A(_02111_),
    .B(_02192_),
    .C(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21o_1 _09293_ (.A1(_02192_),
    .A2(_02193_),
    .B1(_02111_),
    .X(_02195_));
 sky130_fd_sc_hd__and2_1 _09294_ (.A(_02194_),
    .B(_02195_),
    .X(_02197_));
 sky130_fd_sc_hd__nor3_1 _09295_ (.A(_01601_),
    .B(_01691_),
    .C(_01692_),
    .Y(_02198_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(_01593_),
    .B(_01594_),
    .X(_02199_));
 sky130_fd_sc_hd__o21a_1 _09297_ (.A1(_01581_),
    .A2(_01595_),
    .B1(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__nor2_1 _09298_ (.A(_01065_),
    .B(_01624_),
    .Y(_02201_));
 sky130_fd_sc_hd__a31o_1 _09299_ (.A1(_00059_),
    .A2(_00062_),
    .A3(_01556_),
    .B1(_01555_),
    .X(_02202_));
 sky130_fd_sc_hd__a22o_1 _09300_ (.A1(net175),
    .A2(net134),
    .B1(net145),
    .B2(net174),
    .X(_02203_));
 sky130_fd_sc_hd__nand4_2 _09301_ (.A(net174),
    .B(net175),
    .C(_00985_),
    .D(net145),
    .Y(_02204_));
 sky130_fd_sc_hd__a22o_1 _09302_ (.A1(net176),
    .A2(_00479_),
    .B1(_02203_),
    .B2(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__nand4_1 _09303_ (.A(net176),
    .B(_00479_),
    .C(_02203_),
    .D(_02204_),
    .Y(_02206_));
 sky130_fd_sc_hd__and3_1 _09304_ (.A(_01565_),
    .B(_02205_),
    .C(_02206_),
    .X(_02208_));
 sky130_fd_sc_hd__a21o_1 _09305_ (.A1(_02205_),
    .A2(_02206_),
    .B1(_01565_),
    .X(_02209_));
 sky130_fd_sc_hd__or2b_1 _09306_ (.A(_02208_),
    .B_N(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__xor2_1 _09307_ (.A(_02202_),
    .B(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__a22oi_2 _09308_ (.A1(net183),
    .A2(net197),
    .B1(net198),
    .B2(net182),
    .Y(_02212_));
 sky130_fd_sc_hd__and4_1 _09309_ (.A(net183),
    .B(net182),
    .C(net197),
    .D(net198),
    .X(_02213_));
 sky130_fd_sc_hd__nor2_1 _09310_ (.A(_02212_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__buf_2 _09311_ (.A(net156),
    .X(_02215_));
 sky130_fd_sc_hd__nand2_1 _09312_ (.A(net167),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__xnor2_1 _09313_ (.A(_02214_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__and4_1 _09314_ (.A(net184),
    .B(_00049_),
    .C(_00058_),
    .D(_00481_),
    .X(_02219_));
 sky130_fd_sc_hd__and4_1 _09315_ (.A(net183),
    .B(_01567_),
    .C(_01568_),
    .D(_01569_),
    .X(_02220_));
 sky130_fd_sc_hd__a22o_1 _09316_ (.A1(_00989_),
    .A2(net186),
    .B1(net195),
    .B2(net185),
    .X(_02221_));
 sky130_fd_sc_hd__nand4_2 _09317_ (.A(_00047_),
    .B(_00989_),
    .C(net186),
    .D(_00480_),
    .Y(_02222_));
 sky130_fd_sc_hd__a22o_1 _09318_ (.A1(_05115_),
    .A2(_01567_),
    .B1(_02221_),
    .B2(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__nand4_2 _09319_ (.A(_05115_),
    .B(_01567_),
    .C(_02221_),
    .D(_02222_),
    .Y(_02224_));
 sky130_fd_sc_hd__o211ai_2 _09320_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_02223_),
    .C1(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__a211o_1 _09321_ (.A1(_02223_),
    .A2(_02224_),
    .B1(_02219_),
    .C1(_02220_),
    .X(_02226_));
 sky130_fd_sc_hd__nand3_1 _09322_ (.A(_02217_),
    .B(_02225_),
    .C(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__a21o_1 _09323_ (.A1(_02225_),
    .A2(_02226_),
    .B1(_02217_),
    .X(_02228_));
 sky130_fd_sc_hd__a21bo_1 _09324_ (.A1(_01566_),
    .A2(_01574_),
    .B1_N(_01573_),
    .X(_02230_));
 sky130_fd_sc_hd__and3_2 _09325_ (.A(_02227_),
    .B(_02228_),
    .C(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__a21oi_1 _09326_ (.A1(_02227_),
    .A2(_02228_),
    .B1(_02230_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor3_1 _09327_ (.A(_02211_),
    .B(_02231_),
    .C(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__o21a_1 _09328_ (.A1(_02231_),
    .A2(_02232_),
    .B1(_02211_),
    .X(_02234_));
 sky130_fd_sc_hd__and2b_1 _09329_ (.A_N(_01589_),
    .B(_01590_),
    .X(_02235_));
 sky130_fd_sc_hd__a21o_1 _09330_ (.A1(_01606_),
    .A2(_01614_),
    .B1(_01613_),
    .X(_02236_));
 sky130_fd_sc_hd__a32o_1 _09331_ (.A1(_05093_),
    .A2(_00489_),
    .A3(_01586_),
    .B1(_01585_),
    .B2(_01584_),
    .X(_02237_));
 sky130_fd_sc_hd__a22o_1 _09332_ (.A1(net192),
    .A2(net188),
    .B1(net189),
    .B2(net191),
    .X(_02238_));
 sky130_fd_sc_hd__clkbuf_4 _09333_ (.A(net189),
    .X(_02239_));
 sky130_fd_sc_hd__nand4_2 _09334_ (.A(net191),
    .B(net192),
    .C(net188),
    .D(_02239_),
    .Y(_02241_));
 sky130_fd_sc_hd__a22o_1 _09335_ (.A1(_05093_),
    .A2(_01002_),
    .B1(_02238_),
    .B2(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__nand4_2 _09336_ (.A(net193),
    .B(_01002_),
    .C(_02238_),
    .D(_02241_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand3_2 _09337_ (.A(_01605_),
    .B(_02242_),
    .C(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__a21o_1 _09338_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_01605_),
    .X(_02245_));
 sky130_fd_sc_hd__nand3_2 _09339_ (.A(_02237_),
    .B(_02244_),
    .C(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21o_1 _09340_ (.A1(_02244_),
    .A2(_02245_),
    .B1(_02237_),
    .X(_02247_));
 sky130_fd_sc_hd__nand3_1 _09341_ (.A(_02236_),
    .B(_02246_),
    .C(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__a21o_1 _09342_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02236_),
    .X(_02249_));
 sky130_fd_sc_hd__nand3_1 _09343_ (.A(_02235_),
    .B(_02248_),
    .C(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21o_1 _09344_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02235_),
    .X(_02252_));
 sky130_fd_sc_hd__and2b_1 _09345_ (.A_N(_01591_),
    .B(_01583_),
    .X(_02253_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(_01582_),
    .A2(_01592_),
    .B1(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__nand3_2 _09347_ (.A(_02250_),
    .B(_02252_),
    .C(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__a21o_1 _09348_ (.A1(_02250_),
    .A2(_02252_),
    .B1(_02254_),
    .X(_02256_));
 sky130_fd_sc_hd__or4bb_2 _09349_ (.A(_02233_),
    .B(_02234_),
    .C_N(_02255_),
    .D_N(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__a2bb2o_1 _09350_ (.A1_N(_02233_),
    .A2_N(_02234_),
    .B1(_02255_),
    .B2(_02256_),
    .X(_02258_));
 sky130_fd_sc_hd__o211a_1 _09351_ (.A1(_02201_),
    .A2(_01626_),
    .B1(_02257_),
    .C1(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__a211oi_1 _09352_ (.A1(_02257_),
    .A2(_02258_),
    .B1(_02201_),
    .C1(_01626_),
    .Y(_02260_));
 sky130_fd_sc_hd__nor3_1 _09353_ (.A(_02200_),
    .B(_02259_),
    .C(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__o21a_1 _09354_ (.A1(_02259_),
    .A2(_02260_),
    .B1(_02200_),
    .X(_02263_));
 sky130_fd_sc_hd__nor2_2 _09355_ (.A(_02261_),
    .B(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _09356_ (.A(_01616_),
    .B(_01623_),
    .Y(_02265_));
 sky130_fd_sc_hd__a31o_1 _09357_ (.A1(_00513_),
    .A2(_01036_),
    .A3(_01622_),
    .B1(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__or3b_1 _09358_ (.A(_01642_),
    .B(_01643_),
    .C_N(_01069_),
    .X(_02267_));
 sky130_fd_sc_hd__a22oi_2 _09359_ (.A1(net219),
    .A2(net231),
    .B1(net232),
    .B2(net218),
    .Y(_02268_));
 sky130_fd_sc_hd__and4_1 _09360_ (.A(net218),
    .B(net219),
    .C(net231),
    .D(net232),
    .X(_02269_));
 sky130_fd_sc_hd__or2_1 _09361_ (.A(_02268_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__nand2_1 _09362_ (.A(net217),
    .B(net233),
    .Y(_02271_));
 sky130_fd_sc_hd__xnor2_1 _09363_ (.A(_02270_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__a22o_1 _09364_ (.A1(net229),
    .A2(net221),
    .B1(net222),
    .B2(net228),
    .X(_02274_));
 sky130_fd_sc_hd__nand4_1 _09365_ (.A(net228),
    .B(net229),
    .C(net221),
    .D(net222),
    .Y(_02275_));
 sky130_fd_sc_hd__a22oi_2 _09366_ (.A1(_00080_),
    .A2(_00516_),
    .B1(_02274_),
    .B2(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__and4_2 _09367_ (.A(_00080_),
    .B(net230),
    .C(_02274_),
    .D(_02275_),
    .X(_02277_));
 sky130_fd_sc_hd__or2_1 _09368_ (.A(_02276_),
    .B(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(_01610_),
    .B(_01611_),
    .Y(_02279_));
 sky130_fd_sc_hd__xnor2_1 _09370_ (.A(_02278_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__xnor2_1 _09371_ (.A(_02272_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__a32o_1 _09372_ (.A1(net32),
    .A2(net48),
    .A3(_01632_),
    .B1(_01631_),
    .B2(_00530_),
    .X(_02282_));
 sky130_fd_sc_hd__nand4_1 _09373_ (.A(net32),
    .B(net226),
    .C(net49),
    .D(net225),
    .Y(_02283_));
 sky130_fd_sc_hd__a22o_1 _09374_ (.A1(net32),
    .A2(net49),
    .B1(net225),
    .B2(net226),
    .X(_02285_));
 sky130_fd_sc_hd__a22o_1 _09375_ (.A1(net227),
    .A2(net224),
    .B1(_02283_),
    .B2(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__nand4_1 _09376_ (.A(net227),
    .B(net224),
    .C(_02283_),
    .D(_02285_),
    .Y(_02287_));
 sky130_fd_sc_hd__and3_1 _09377_ (.A(_02282_),
    .B(_02286_),
    .C(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__a21oi_1 _09378_ (.A1(_02286_),
    .A2(_02287_),
    .B1(_02282_),
    .Y(_02289_));
 sky130_fd_sc_hd__or3_1 _09379_ (.A(_01619_),
    .B(_02288_),
    .C(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__o21ai_1 _09380_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_01619_),
    .Y(_02291_));
 sky130_fd_sc_hd__o21a_1 _09381_ (.A1(_01038_),
    .A2(_01620_),
    .B1(_01621_),
    .X(_02292_));
 sky130_fd_sc_hd__nand3_1 _09382_ (.A(_02290_),
    .B(_02291_),
    .C(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__a21o_1 _09383_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02292_),
    .X(_02294_));
 sky130_fd_sc_hd__and3_1 _09384_ (.A(_02281_),
    .B(_02293_),
    .C(_02294_),
    .X(_02296_));
 sky130_fd_sc_hd__a21oi_1 _09385_ (.A1(_02293_),
    .A2(_02294_),
    .B1(_02281_),
    .Y(_02297_));
 sky130_fd_sc_hd__a211o_1 _09386_ (.A1(_02267_),
    .A2(_01646_),
    .B1(_02296_),
    .C1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__o211ai_2 _09387_ (.A1(_02296_),
    .A2(_02297_),
    .B1(_02267_),
    .C1(_01646_),
    .Y(_02299_));
 sky130_fd_sc_hd__and3_1 _09388_ (.A(_02266_),
    .B(_02298_),
    .C(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__a21oi_1 _09389_ (.A1(_02298_),
    .A2(_02299_),
    .B1(_02266_),
    .Y(_02301_));
 sky130_fd_sc_hd__nor2_2 _09390_ (.A(_02300_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__a21boi_2 _09391_ (.A1(_01634_),
    .A2(_01641_),
    .B1_N(_01640_),
    .Y(_02303_));
 sky130_fd_sc_hd__a22oi_2 _09392_ (.A1(net36),
    .A2(_00530_),
    .B1(_01051_),
    .B2(_04906_),
    .Y(_02304_));
 sky130_fd_sc_hd__and4_1 _09393_ (.A(_04906_),
    .B(net36),
    .C(net46),
    .D(net47),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_1 _09394_ (.A(_02304_),
    .B(_02305_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(_03084_),
    .B(net48),
    .Y(_02308_));
 sky130_fd_sc_hd__xnor2_1 _09396_ (.A(_02307_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__and4_1 _09397_ (.A(_03194_),
    .B(_04862_),
    .C(_00543_),
    .D(_01068_),
    .X(_02310_));
 sky130_fd_sc_hd__and4_1 _09398_ (.A(_00107_),
    .B(_00097_),
    .C(_01635_),
    .D(_01636_),
    .X(_02311_));
 sky130_fd_sc_hd__a22o_1 _09399_ (.A1(net43),
    .A2(net38),
    .B1(net39),
    .B2(net42),
    .X(_02312_));
 sky130_fd_sc_hd__nand4_1 _09400_ (.A(_03194_),
    .B(net43),
    .C(_01068_),
    .D(net39),
    .Y(_02313_));
 sky130_fd_sc_hd__and2_1 _09401_ (.A(net44),
    .B(net37),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _09402_ (.A1(_02312_),
    .A2(_02313_),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__nand3_1 _09403_ (.A(_02312_),
    .B(_02313_),
    .C(_02314_),
    .Y(_02316_));
 sky130_fd_sc_hd__o211ai_2 _09404_ (.A1(_02310_),
    .A2(_02311_),
    .B1(_02315_),
    .C1(_02316_),
    .Y(_02318_));
 sky130_fd_sc_hd__a211o_1 _09405_ (.A1(_02315_),
    .A2(_02316_),
    .B1(_02310_),
    .C1(_02311_),
    .X(_02319_));
 sky130_fd_sc_hd__nand3_1 _09406_ (.A(_02309_),
    .B(_02318_),
    .C(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__a21o_1 _09407_ (.A1(_02318_),
    .A2(_02319_),
    .B1(_02309_),
    .X(_02321_));
 sky130_fd_sc_hd__and3_1 _09408_ (.A(_01657_),
    .B(_02320_),
    .C(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__a21oi_1 _09409_ (.A1(_02320_),
    .A2(_02321_),
    .B1(_01657_),
    .Y(_02323_));
 sky130_fd_sc_hd__nor2_1 _09410_ (.A(_02322_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_2 _09411_ (.A(_02303_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__inv_2 _09412_ (.A(_01678_),
    .Y(_02326_));
 sky130_fd_sc_hd__a31o_1 _09413_ (.A1(_03095_),
    .A2(_01072_),
    .A3(_01662_),
    .B1(_01661_),
    .X(_02327_));
 sky130_fd_sc_hd__clkbuf_4 _09414_ (.A(net40),
    .X(_02329_));
 sky130_fd_sc_hd__a22o_1 _09415_ (.A1(_03095_),
    .A2(net56),
    .B1(net67),
    .B2(net1),
    .X(_02330_));
 sky130_fd_sc_hd__nand4_2 _09416_ (.A(_03095_),
    .B(net1),
    .C(net56),
    .D(net67),
    .Y(_02331_));
 sky130_fd_sc_hd__a22o_1 _09417_ (.A1(net41),
    .A2(_02329_),
    .B1(_02330_),
    .B2(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__nand4_1 _09418_ (.A(net41),
    .B(_02329_),
    .C(_02330_),
    .D(_02331_),
    .Y(_02333_));
 sky130_fd_sc_hd__and3_1 _09419_ (.A(_02327_),
    .B(_02332_),
    .C(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__a21o_1 _09420_ (.A1(_02332_),
    .A2(_02333_),
    .B1(_02327_),
    .X(_02335_));
 sky130_fd_sc_hd__and2b_1 _09421_ (.A_N(_02334_),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__xnor2_2 _09422_ (.A(_01655_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__and4_1 _09423_ (.A(net190),
    .B(net23),
    .C(_00550_),
    .D(net34),
    .X(_02338_));
 sky130_fd_sc_hd__a22o_1 _09424_ (.A1(_00109_),
    .A2(_00550_),
    .B1(_00544_),
    .B2(_00549_),
    .X(_02340_));
 sky130_fd_sc_hd__and2b_1 _09425_ (.A_N(_02338_),
    .B(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__nand2_1 _09426_ (.A(_04939_),
    .B(_01072_),
    .Y(_02342_));
 sky130_fd_sc_hd__xnor2_1 _09427_ (.A(_02341_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__and2_1 _09428_ (.A(net12),
    .B(_01666_),
    .X(_02344_));
 sky130_fd_sc_hd__nand4_1 _09429_ (.A(_02789_),
    .B(_03106_),
    .C(net223),
    .D(net234),
    .Y(_02345_));
 sky130_fd_sc_hd__a22o_1 _09430_ (.A1(_03106_),
    .A2(net223),
    .B1(net234),
    .B2(_02789_),
    .X(_02346_));
 sky130_fd_sc_hd__nand3_1 _09431_ (.A(_02344_),
    .B(_02345_),
    .C(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a21o_1 _09432_ (.A1(_02345_),
    .A2(_02346_),
    .B1(_02344_),
    .X(_02348_));
 sky130_fd_sc_hd__a21bo_1 _09433_ (.A1(_01665_),
    .A2(_01669_),
    .B1_N(_01668_),
    .X(_02349_));
 sky130_fd_sc_hd__nand3_1 _09434_ (.A(_02347_),
    .B(_02348_),
    .C(_02349_),
    .Y(_02351_));
 sky130_fd_sc_hd__a21o_1 _09435_ (.A1(_02347_),
    .A2(_02348_),
    .B1(_02349_),
    .X(_02352_));
 sky130_fd_sc_hd__nand3_1 _09436_ (.A(_02343_),
    .B(_02351_),
    .C(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21o_1 _09437_ (.A1(_02351_),
    .A2(_02352_),
    .B1(_02343_),
    .X(_02354_));
 sky130_fd_sc_hd__a21bo_1 _09438_ (.A1(_01664_),
    .A2(_01674_),
    .B1_N(_01673_),
    .X(_02355_));
 sky130_fd_sc_hd__and3_1 _09439_ (.A(_02353_),
    .B(_02354_),
    .C(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_2 _09440_ (.A1(_02353_),
    .A2(_02354_),
    .B1(_02355_),
    .Y(_02357_));
 sky130_fd_sc_hd__or3_2 _09441_ (.A(_02337_),
    .B(_02356_),
    .C(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__o21ai_2 _09442_ (.A1(_02356_),
    .A2(_02357_),
    .B1(_02337_),
    .Y(_02359_));
 sky130_fd_sc_hd__o211ai_2 _09443_ (.A1(_02326_),
    .A2(_01680_),
    .B1(_02358_),
    .C1(_02359_),
    .Y(_02360_));
 sky130_fd_sc_hd__a211o_2 _09444_ (.A1(_02358_),
    .A2(_02359_),
    .B1(_02326_),
    .C1(_01680_),
    .X(_02362_));
 sky130_fd_sc_hd__and3_2 _09445_ (.A(_02325_),
    .B(_02360_),
    .C(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__a21oi_2 _09446_ (.A1(_02360_),
    .A2(_02362_),
    .B1(_02325_),
    .Y(_02364_));
 sky130_fd_sc_hd__a211o_1 _09447_ (.A1(_01682_),
    .A2(_01684_),
    .B1(_02363_),
    .C1(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__o211ai_4 _09448_ (.A1(_02363_),
    .A2(_02364_),
    .B1(_01682_),
    .C1(_01684_),
    .Y(_02366_));
 sky130_fd_sc_hd__and3_2 _09449_ (.A(_02302_),
    .B(_02365_),
    .C(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a21oi_2 _09450_ (.A1(_02365_),
    .A2(_02366_),
    .B1(_02302_),
    .Y(_02368_));
 sky130_fd_sc_hd__a211o_1 _09451_ (.A1(_01686_),
    .A2(_01688_),
    .B1(_02367_),
    .C1(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__o211ai_4 _09452_ (.A1(_02367_),
    .A2(_02368_),
    .B1(_01686_),
    .C1(net311),
    .Y(_02370_));
 sky130_fd_sc_hd__nand3_1 _09453_ (.A(_02264_),
    .B(_02369_),
    .C(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__a21o_1 _09454_ (.A1(_02369_),
    .A2(_02370_),
    .B1(_02264_),
    .X(_02373_));
 sky130_fd_sc_hd__o211ai_2 _09455_ (.A1(_01691_),
    .A2(_02198_),
    .B1(_02371_),
    .C1(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a211o_1 _09456_ (.A1(_02371_),
    .A2(_02373_),
    .B1(_01691_),
    .C1(_02198_),
    .X(_02375_));
 sky130_fd_sc_hd__nand3_1 _09457_ (.A(_02197_),
    .B(_02374_),
    .C(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _09458_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02197_),
    .X(_02377_));
 sky130_fd_sc_hd__o211ai_2 _09459_ (.A1(_01695_),
    .A2(_02110_),
    .B1(_02376_),
    .C1(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a211o_1 _09460_ (.A1(_02376_),
    .A2(_02377_),
    .B1(_01695_),
    .C1(_02110_),
    .X(_02379_));
 sky130_fd_sc_hd__nand3_1 _09461_ (.A(_02109_),
    .B(_02378_),
    .C(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__a21o_1 _09462_ (.A1(_02378_),
    .A2(_02379_),
    .B1(_02109_),
    .X(_02381_));
 sky130_fd_sc_hd__o211ai_2 _09463_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_02380_),
    .C1(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__a211o_1 _09464_ (.A1(_02380_),
    .A2(_02381_),
    .B1(_01974_),
    .C1(_01975_),
    .X(_02384_));
 sky130_fd_sc_hd__nand3_1 _09465_ (.A(_01973_),
    .B(_02382_),
    .C(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__a21o_1 _09466_ (.A1(_02382_),
    .A2(_02384_),
    .B1(_01973_),
    .X(_02386_));
 sky130_fd_sc_hd__o211ai_2 _09467_ (.A1(_01765_),
    .A2(_01766_),
    .B1(_02385_),
    .C1(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__a211o_1 _09468_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_01765_),
    .C1(_01766_),
    .X(_02388_));
 sky130_fd_sc_hd__nand3_2 _09469_ (.A(_01764_),
    .B(_02387_),
    .C(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__a21o_1 _09470_ (.A1(_02387_),
    .A2(_02388_),
    .B1(_01764_),
    .X(_02390_));
 sky130_fd_sc_hd__o211ai_4 _09471_ (.A1(_01728_),
    .A2(_01710_),
    .B1(_02389_),
    .C1(_02390_),
    .Y(_02391_));
 sky130_fd_sc_hd__a211o_1 _09472_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_01728_),
    .C1(_01710_),
    .X(_02392_));
 sky130_fd_sc_hd__nand3_2 _09473_ (.A(_01727_),
    .B(_02391_),
    .C(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__a21o_1 _09474_ (.A1(_02391_),
    .A2(_02392_),
    .B1(_01727_),
    .X(_02395_));
 sky130_fd_sc_hd__o211a_1 _09475_ (.A1(_01712_),
    .A2(net286),
    .B1(_02393_),
    .C1(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__a211oi_1 _09476_ (.A1(_02393_),
    .A2(_02395_),
    .B1(_01712_),
    .C1(net286),
    .Y(_02397_));
 sky130_fd_sc_hd__nor2_1 _09477_ (.A(_02396_),
    .B(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__and2b_1 _09478_ (.A_N(_01716_),
    .B(_01717_),
    .X(_02399_));
 sky130_fd_sc_hd__a31o_1 _09479_ (.A1(_01132_),
    .A2(_01133_),
    .A3(_01718_),
    .B1(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__xor2_1 _09480_ (.A(_02398_),
    .B(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__and2_1 _09481_ (.A(net283),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__or2_1 _09482_ (.A(net283),
    .B(_02401_),
    .X(_02403_));
 sky130_fd_sc_hd__or2b_1 _09483_ (.A(_02402_),
    .B_N(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__a21o_1 _09484_ (.A1(_01721_),
    .A2(_01724_),
    .B1(_01720_),
    .X(_02406_));
 sky130_fd_sc_hd__xor2_1 _09485_ (.A(_02404_),
    .B(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__nor2_1 _09486_ (.A(_00166_),
    .B(_02407_),
    .Y(_00007_));
 sky130_fd_sc_hd__or2b_1 _09487_ (.A(_01763_),
    .B_N(_01729_),
    .X(_02408_));
 sky130_fd_sc_hd__o21ai_1 _09488_ (.A1(_01730_),
    .A2(_01762_),
    .B1(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__or2b_1 _09489_ (.A(_01733_),
    .B_N(_01760_),
    .X(_02410_));
 sky130_fd_sc_hd__a21bo_1 _09490_ (.A1(_01731_),
    .A2(_01761_),
    .B1_N(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__and2_2 _09491_ (.A(_01969_),
    .B(_01971_),
    .X(_02412_));
 sky130_fd_sc_hd__and2_1 _09492_ (.A(_01159_),
    .B(_01160_),
    .X(_02413_));
 sky130_fd_sc_hd__a32o_2 _09493_ (.A1(_01735_),
    .A2(_01756_),
    .A3(_01757_),
    .B1(_01759_),
    .B2(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__nand2_4 _09494_ (.A(_01894_),
    .B(_01896_),
    .Y(_02416_));
 sky130_fd_sc_hd__o21ai_4 _09495_ (.A1(_01751_),
    .A2(_01752_),
    .B1(_01757_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_2 _09496_ (.A(_01799_),
    .B(_01801_),
    .Y(_02418_));
 sky130_fd_sc_hd__or2_1 _09497_ (.A(_01780_),
    .B(_01782_),
    .X(_02419_));
 sky130_fd_sc_hd__a22o_1 _09498_ (.A1(net161),
    .A2(net170),
    .B1(net162),
    .B2(net169),
    .X(_02420_));
 sky130_fd_sc_hd__nand4_1 _09499_ (.A(net169),
    .B(net161),
    .C(_00171_),
    .D(_01777_),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(_02420_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _09501_ (.A(_06243_),
    .B(net171),
    .Y(_02423_));
 sky130_fd_sc_hd__xnor2_1 _09502_ (.A(_02422_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__xnor2_1 _09503_ (.A(_02419_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__o21ba_1 _09504_ (.A1(_01737_),
    .A2(_01740_),
    .B1_N(_01738_),
    .X(_02427_));
 sky130_fd_sc_hd__xor2_1 _09505_ (.A(_02425_),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__and2b_1 _09506_ (.A_N(_01736_),
    .B(_01741_),
    .X(_02429_));
 sky130_fd_sc_hd__a21oi_1 _09507_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__or2_1 _09508_ (.A(_02428_),
    .B(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__nand2_1 _09509_ (.A(_02428_),
    .B(_02430_),
    .Y(_02432_));
 sky130_fd_sc_hd__and2_1 _09510_ (.A(_02431_),
    .B(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__and2_1 _09511_ (.A(_06127_),
    .B(_01157_),
    .X(_02434_));
 sky130_fd_sc_hd__or2_1 _09512_ (.A(_02433_),
    .B(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(_02433_),
    .B(_02434_),
    .Y(_02436_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(_02435_),
    .B(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__o21ba_1 _09515_ (.A1(_01744_),
    .A2(_01746_),
    .B1_N(_01750_),
    .X(_02439_));
 sky130_fd_sc_hd__xor2_1 _09516_ (.A(_02438_),
    .B(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__and2_1 _09517_ (.A(_04227_),
    .B(net173),
    .X(_02441_));
 sky130_fd_sc_hd__nor2_1 _09518_ (.A(_02440_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__and2_1 _09519_ (.A(_02440_),
    .B(_02441_),
    .X(_02443_));
 sky130_fd_sc_hd__or2_2 _09520_ (.A(_02442_),
    .B(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__xor2_4 _09521_ (.A(_02418_),
    .B(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__xor2_4 _09522_ (.A(_02417_),
    .B(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__xnor2_4 _09523_ (.A(_02416_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__xnor2_4 _09524_ (.A(_02414_),
    .B(_02447_),
    .Y(_02449_));
 sky130_fd_sc_hd__xnor2_2 _09525_ (.A(_02412_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__xnor2_2 _09526_ (.A(_02411_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__o211a_1 _09527_ (.A1(_01345_),
    .A2(_01898_),
    .B1(_01963_),
    .C1(_01964_),
    .X(_02452_));
 sky130_fd_sc_hd__or2_2 _09528_ (.A(_02452_),
    .B(_01967_),
    .X(_02453_));
 sky130_fd_sc_hd__and2_2 _09529_ (.A(_01795_),
    .B(_01797_),
    .X(_02454_));
 sky130_fd_sc_hd__or2_2 _09530_ (.A(_01817_),
    .B(_01849_),
    .X(_02455_));
 sky130_fd_sc_hd__and2b_1 _09531_ (.A_N(_01776_),
    .B(_01792_),
    .X(_02456_));
 sky130_fd_sc_hd__a21o_2 _09532_ (.A1(_01775_),
    .A2(_01793_),
    .B1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_2 _09533_ (.A(_01844_),
    .B(_01846_),
    .Y(_02458_));
 sky130_fd_sc_hd__or2_1 _09534_ (.A(_01184_),
    .B(_01790_),
    .X(_02460_));
 sky130_fd_sc_hd__o31ai_4 _09535_ (.A1(_01781_),
    .A2(_01782_),
    .A3(_01791_),
    .B1(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__or2b_1 _09536_ (.A(_01825_),
    .B_N(_01819_),
    .X(_02462_));
 sky130_fd_sc_hd__a21bo_2 _09537_ (.A1(_01220_),
    .A2(_01824_),
    .B1_N(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_4 _09538_ (.A(net164),
    .X(_02464_));
 sky130_fd_sc_hd__a22oi_1 _09539_ (.A1(_06130_),
    .A2(_01188_),
    .B1(_02464_),
    .B2(_04238_),
    .Y(_02465_));
 sky130_fd_sc_hd__and4_1 _09540_ (.A(_04238_),
    .B(_06130_),
    .C(_01188_),
    .D(net164),
    .X(_02466_));
 sky130_fd_sc_hd__or2_2 _09541_ (.A(_02465_),
    .B(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__a22o_1 _09542_ (.A1(net18),
    .A2(net29),
    .B1(net30),
    .B2(net17),
    .X(_02468_));
 sky130_fd_sc_hd__inv_2 _09543_ (.A(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__and4_1 _09544_ (.A(net17),
    .B(net18),
    .C(net29),
    .D(net30),
    .X(_02471_));
 sky130_fd_sc_hd__o2bb2a_1 _09545_ (.A1_N(_04435_),
    .A2_N(_01784_),
    .B1(_02469_),
    .B2(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__and4b_1 _09546_ (.A_N(_02471_),
    .B(net31),
    .C(_04435_),
    .D(_02468_),
    .X(_02473_));
 sky130_fd_sc_hd__or2_2 _09547_ (.A(_02472_),
    .B(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__nor2_1 _09548_ (.A(_01787_),
    .B(_01789_),
    .Y(_02475_));
 sky130_fd_sc_hd__xnor2_2 _09549_ (.A(_02474_),
    .B(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__xnor2_2 _09550_ (.A(_02467_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__xor2_4 _09551_ (.A(_02463_),
    .B(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__xor2_4 _09552_ (.A(_02461_),
    .B(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__xnor2_4 _09553_ (.A(_02458_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__xnor2_4 _09554_ (.A(_02457_),
    .B(_02480_),
    .Y(_02482_));
 sky130_fd_sc_hd__xnor2_4 _09555_ (.A(_02455_),
    .B(_02482_),
    .Y(_02483_));
 sky130_fd_sc_hd__xnor2_4 _09556_ (.A(_02454_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _09557_ (.A(_01821_),
    .B(_01823_),
    .Y(_02485_));
 sky130_fd_sc_hd__a21bo_1 _09558_ (.A1(_01829_),
    .A2(_01831_),
    .B1_N(_01830_),
    .X(_02486_));
 sky130_fd_sc_hd__a22o_1 _09559_ (.A1(net27),
    .A2(net20),
    .B1(net21),
    .B2(net26),
    .X(_02487_));
 sky130_fd_sc_hd__nand4_2 _09560_ (.A(_06142_),
    .B(_06264_),
    .C(net20),
    .D(_01217_),
    .Y(_02488_));
 sky130_fd_sc_hd__a22o_1 _09561_ (.A1(_00239_),
    .A2(net28),
    .B1(_02487_),
    .B2(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__nand4_2 _09562_ (.A(_00239_),
    .B(_00250_),
    .C(_02487_),
    .D(_02488_),
    .Y(_02490_));
 sky130_fd_sc_hd__and3_1 _09563_ (.A(_02486_),
    .B(_02489_),
    .C(_02490_),
    .X(_02491_));
 sky130_fd_sc_hd__a21oi_1 _09564_ (.A1(_02489_),
    .A2(_02490_),
    .B1(_02486_),
    .Y(_02493_));
 sky130_fd_sc_hd__nor2_1 _09565_ (.A(_02491_),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__xnor2_1 _09566_ (.A(_02485_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(_01840_),
    .B(_01841_),
    .Y(_02496_));
 sky130_fd_sc_hd__or2_1 _09568_ (.A(_01834_),
    .B(_01842_),
    .X(_02497_));
 sky130_fd_sc_hd__buf_2 _09569_ (.A(net22),
    .X(_02498_));
 sky130_fd_sc_hd__a22oi_2 _09570_ (.A1(_04292_),
    .A2(net102),
    .B1(_02498_),
    .B2(_04446_),
    .Y(_02499_));
 sky130_fd_sc_hd__and4_2 _09571_ (.A(_04292_),
    .B(_04446_),
    .C(net102),
    .D(_02498_),
    .X(_02500_));
 sky130_fd_sc_hd__nor2_1 _09572_ (.A(_02499_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__a22o_1 _09573_ (.A1(_00200_),
    .A2(_00238_),
    .B1(_00703_),
    .B2(net88),
    .X(_02502_));
 sky130_fd_sc_hd__nand4_1 _09574_ (.A(_06284_),
    .B(_00200_),
    .C(_00238_),
    .D(_00703_),
    .Y(_02504_));
 sky130_fd_sc_hd__a22o_1 _09575_ (.A1(_06159_),
    .A2(_01835_),
    .B1(_02502_),
    .B2(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__nand4_1 _09576_ (.A(_06159_),
    .B(_01835_),
    .C(_02502_),
    .D(_02504_),
    .Y(_02506_));
 sky130_fd_sc_hd__o211a_1 _09577_ (.A1(_01837_),
    .A2(_01839_),
    .B1(_02505_),
    .C1(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a211oi_1 _09578_ (.A1(_02505_),
    .A2(_02506_),
    .B1(_01837_),
    .C1(_01839_),
    .Y(_02508_));
 sky130_fd_sc_hd__or2_1 _09579_ (.A(_02507_),
    .B(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__xor2_1 _09580_ (.A(_02501_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__a21o_1 _09581_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__nand3_1 _09582_ (.A(_02496_),
    .B(_02497_),
    .C(_02510_),
    .Y(_02512_));
 sky130_fd_sc_hd__nand3_1 _09583_ (.A(_02495_),
    .B(_02511_),
    .C(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__a21o_1 _09584_ (.A1(_02511_),
    .A2(_02512_),
    .B1(_02495_),
    .X(_02515_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(_02513_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__and2b_1 _09586_ (.A_N(_01806_),
    .B(_01814_),
    .X(_02517_));
 sky130_fd_sc_hd__and2_1 _09587_ (.A(_01234_),
    .B(_01815_),
    .X(_02518_));
 sky130_fd_sc_hd__and2b_1 _09588_ (.A_N(_01813_),
    .B(_01807_),
    .X(_02519_));
 sky130_fd_sc_hd__a21oi_1 _09589_ (.A1(_01253_),
    .A2(_01812_),
    .B1(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21boi_1 _09590_ (.A1(_01860_),
    .A2(_01867_),
    .B1_N(_01866_),
    .Y(_02521_));
 sky130_fd_sc_hd__a41o_1 _09591_ (.A1(_04424_),
    .A2(_06134_),
    .A3(_00672_),
    .A4(_01251_),
    .B1(_01811_),
    .X(_02522_));
 sky130_fd_sc_hd__o21bai_1 _09592_ (.A1(_01855_),
    .A2(_01859_),
    .B1_N(_01856_),
    .Y(_02523_));
 sky130_fd_sc_hd__a22o_1 _09593_ (.A1(_06254_),
    .A2(net92),
    .B1(_01858_),
    .B2(_04413_),
    .X(_02524_));
 sky130_fd_sc_hd__nand4_2 _09594_ (.A(_04413_),
    .B(_06254_),
    .C(net92),
    .D(_01858_),
    .Y(_02526_));
 sky130_fd_sc_hd__a22o_1 _09595_ (.A1(_06253_),
    .A2(_00672_),
    .B1(_02524_),
    .B2(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__nand4_2 _09596_ (.A(net97),
    .B(_00672_),
    .C(_02524_),
    .D(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand3_1 _09597_ (.A(_02523_),
    .B(_02527_),
    .C(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__a21o_1 _09598_ (.A1(_02527_),
    .A2(_02528_),
    .B1(_02523_),
    .X(_02530_));
 sky130_fd_sc_hd__nand2_1 _09599_ (.A(_02529_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__xor2_1 _09600_ (.A(_02522_),
    .B(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__nor2_1 _09601_ (.A(_02521_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__and2_1 _09602_ (.A(_02521_),
    .B(_02532_),
    .X(_02534_));
 sky130_fd_sc_hd__or3_1 _09603_ (.A(_02520_),
    .B(_02533_),
    .C(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__o21ai_1 _09604_ (.A1(_02533_),
    .A2(_02534_),
    .B1(_02520_),
    .Y(_02537_));
 sky130_fd_sc_hd__o211a_1 _09605_ (.A1(_02517_),
    .A2(_02518_),
    .B1(_02535_),
    .C1(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__a211oi_1 _09606_ (.A1(_02535_),
    .A2(_02537_),
    .B1(_02517_),
    .C1(_02518_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor3_1 _09607_ (.A(_02516_),
    .B(_02538_),
    .C(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21a_1 _09608_ (.A1(_02538_),
    .A2(_02539_),
    .B1(_02516_),
    .X(_02541_));
 sky130_fd_sc_hd__nor2_2 _09609_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__a31o_2 _09610_ (.A1(_01871_),
    .A2(_01880_),
    .A3(_01881_),
    .B1(_01884_),
    .X(_02543_));
 sky130_fd_sc_hd__a21o_2 _09611_ (.A1(_01936_),
    .A2(_01952_),
    .B1(_01951_),
    .X(_02544_));
 sky130_fd_sc_hd__a22oi_1 _09612_ (.A1(_06152_),
    .A2(net137),
    .B1(net138),
    .B2(_04303_),
    .Y(_02545_));
 sky130_fd_sc_hd__and4_1 _09613_ (.A(_04303_),
    .B(net124),
    .C(net137),
    .D(net138),
    .X(_02546_));
 sky130_fd_sc_hd__nor2_1 _09614_ (.A(_02545_),
    .B(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__and4_1 _09615_ (.A(net125),
    .B(_06283_),
    .C(_00210_),
    .D(_00201_),
    .X(_02549_));
 sky130_fd_sc_hd__and4_1 _09616_ (.A(net124),
    .B(_00665_),
    .C(_01861_),
    .D(_01862_),
    .X(_02550_));
 sky130_fd_sc_hd__a22o_1 _09617_ (.A1(net126),
    .A2(net135),
    .B1(net127),
    .B2(net133),
    .X(_02551_));
 sky130_fd_sc_hd__nand4_1 _09618_ (.A(_06283_),
    .B(net126),
    .C(_00201_),
    .D(net127),
    .Y(_02552_));
 sky130_fd_sc_hd__a22o_1 _09619_ (.A1(net125),
    .A2(_00665_),
    .B1(_02551_),
    .B2(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__nand4_1 _09620_ (.A(_06274_),
    .B(_00665_),
    .C(_02551_),
    .D(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__o211a_1 _09621_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02553_),
    .C1(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a211o_1 _09622_ (.A1(_02553_),
    .A2(_02554_),
    .B1(_02549_),
    .C1(_02550_),
    .X(_02556_));
 sky130_fd_sc_hd__and2b_1 _09623_ (.A_N(_02555_),
    .B(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__xnor2_2 _09624_ (.A(_02548_),
    .B(_02557_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _09625_ (.A(_01874_),
    .B(_01876_),
    .Y(_02560_));
 sky130_fd_sc_hd__o21bai_2 _09626_ (.A1(_01938_),
    .A2(_01941_),
    .B1_N(_01939_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(net131),
    .B(net129),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(net132),
    .B(net128),
    .Y(_02563_));
 sky130_fd_sc_hd__xor2_1 _09629_ (.A(_02562_),
    .B(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__xor2_1 _09630_ (.A(_02561_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__xor2_1 _09631_ (.A(_02560_),
    .B(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__a21boi_1 _09632_ (.A1(_01878_),
    .A2(_01879_),
    .B1_N(_01877_),
    .Y(_02567_));
 sky130_fd_sc_hd__xnor2_1 _09633_ (.A(_02566_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__xnor2_2 _09634_ (.A(_02559_),
    .B(_02568_),
    .Y(_02570_));
 sky130_fd_sc_hd__xor2_4 _09635_ (.A(_02544_),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__xor2_4 _09636_ (.A(_02543_),
    .B(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__nor2_2 _09637_ (.A(_01886_),
    .B(_01888_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_4 _09638_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__xnor2_4 _09639_ (.A(_02542_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_2 _09640_ (.A(_01890_),
    .B(_01892_),
    .Y(_02576_));
 sky130_fd_sc_hd__xor2_4 _09641_ (.A(_02575_),
    .B(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__xnor2_4 _09642_ (.A(_02484_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__nor3_1 _09643_ (.A(_01899_),
    .B(_01961_),
    .C(_01962_),
    .Y(_02579_));
 sky130_fd_sc_hd__or2_1 _09644_ (.A(_01957_),
    .B(_01959_),
    .X(_02581_));
 sky130_fd_sc_hd__or2b_1 _09645_ (.A(_02053_),
    .B_N(_02052_),
    .X(_02582_));
 sky130_fd_sc_hd__or2b_1 _09646_ (.A(_02003_),
    .B_N(_02054_),
    .X(_02583_));
 sky130_fd_sc_hd__nor2_1 _09647_ (.A(_01934_),
    .B(_01955_),
    .Y(_02584_));
 sky130_fd_sc_hd__nor3_2 _09648_ (.A(_01981_),
    .B(_02000_),
    .C(_02001_),
    .Y(_02585_));
 sky130_fd_sc_hd__and2_1 _09649_ (.A(_01947_),
    .B(_01949_),
    .X(_02586_));
 sky130_fd_sc_hd__a21o_1 _09650_ (.A1(_01311_),
    .A2(_01909_),
    .B1(_01908_),
    .X(_02587_));
 sky130_fd_sc_hd__and3_1 _09651_ (.A(_06177_),
    .B(net142),
    .C(_01288_),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _09652_ (.A1(net142),
    .A2(net153),
    .B1(net154),
    .B2(_06177_),
    .X(_02589_));
 sky130_fd_sc_hd__a21bo_1 _09653_ (.A1(_00749_),
    .A2(_02588_),
    .B1_N(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__clkbuf_4 _09654_ (.A(net155),
    .X(_02592_));
 sky130_fd_sc_hd__nand2_1 _09655_ (.A(_04128_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__xor2_1 _09656_ (.A(_02590_),
    .B(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__inv_2 _09657_ (.A(_01944_),
    .Y(_02595_));
 sky130_fd_sc_hd__a22o_1 _09658_ (.A1(net151),
    .A2(_00774_),
    .B1(net146),
    .B2(net150),
    .X(_02596_));
 sky130_fd_sc_hd__nand4_1 _09659_ (.A(_06171_),
    .B(_06319_),
    .C(_00774_),
    .D(net146),
    .Y(_02597_));
 sky130_fd_sc_hd__and2_1 _09660_ (.A(_00291_),
    .B(_01293_),
    .X(_02598_));
 sky130_fd_sc_hd__a21o_1 _09661_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__nand3_1 _09662_ (.A(_02596_),
    .B(_02597_),
    .C(_02598_),
    .Y(_02600_));
 sky130_fd_sc_hd__o211ai_2 _09663_ (.A1(_02595_),
    .A2(_01946_),
    .B1(_02599_),
    .C1(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__a211o_1 _09664_ (.A1(_02599_),
    .A2(_02600_),
    .B1(_02595_),
    .C1(_01946_),
    .X(_02603_));
 sky130_fd_sc_hd__nand3_1 _09665_ (.A(_02594_),
    .B(_02601_),
    .C(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__a21o_1 _09666_ (.A1(_02601_),
    .A2(_02603_),
    .B1(_02594_),
    .X(_02605_));
 sky130_fd_sc_hd__and3_1 _09667_ (.A(_02587_),
    .B(_02604_),
    .C(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__a21o_1 _09668_ (.A1(_02604_),
    .A2(_02605_),
    .B1(_02587_),
    .X(_02607_));
 sky130_fd_sc_hd__inv_2 _09669_ (.A(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__nor3_1 _09670_ (.A(_02586_),
    .B(_02606_),
    .C(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__o21a_1 _09671_ (.A1(_02606_),
    .A2(_02608_),
    .B1(_02586_),
    .X(_02610_));
 sky130_fd_sc_hd__nand3_1 _09672_ (.A(_01927_),
    .B(_01928_),
    .C(_01929_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_1 _09673_ (.A(_01904_),
    .B(_01907_),
    .Y(_02612_));
 sky130_fd_sc_hd__and4_1 _09674_ (.A(_06086_),
    .B(_06362_),
    .C(_00297_),
    .D(_00757_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_4 _09675_ (.A(net147),
    .X(_02615_));
 sky130_fd_sc_hd__nand4_2 _09676_ (.A(_03941_),
    .B(_04139_),
    .C(net216),
    .D(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__a22o_1 _09677_ (.A1(_03941_),
    .A2(net216),
    .B1(_02615_),
    .B2(_04139_),
    .X(_02617_));
 sky130_fd_sc_hd__o211a_1 _09678_ (.A1(_02614_),
    .A2(_01916_),
    .B1(_02616_),
    .C1(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a211o_1 _09679_ (.A1(_02616_),
    .A2(_02617_),
    .B1(_02614_),
    .C1(_01916_),
    .X(_02619_));
 sky130_fd_sc_hd__and2b_1 _09680_ (.A_N(_02618_),
    .B(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__xnor2_1 _09681_ (.A(_02612_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__and3_1 _09682_ (.A(_06361_),
    .B(_00343_),
    .C(net214),
    .X(_02622_));
 sky130_fd_sc_hd__a22o_1 _09683_ (.A1(net204),
    .A2(net213),
    .B1(net214),
    .B2(_06361_),
    .X(_02623_));
 sky130_fd_sc_hd__a21bo_1 _09684_ (.A1(_00297_),
    .A2(_02622_),
    .B1_N(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__buf_2 _09685_ (.A(net215),
    .X(_02626_));
 sky130_fd_sc_hd__nand2_1 _09686_ (.A(_06086_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__xor2_2 _09687_ (.A(_02625_),
    .B(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__a22o_1 _09688_ (.A1(_06173_),
    .A2(net206),
    .B1(net207),
    .B2(_04106_),
    .X(_02629_));
 sky130_fd_sc_hd__nand4_2 _09689_ (.A(_04106_),
    .B(_06173_),
    .C(net206),
    .D(net207),
    .Y(_02630_));
 sky130_fd_sc_hd__and2_1 _09690_ (.A(net211),
    .B(net205),
    .X(_02631_));
 sky130_fd_sc_hd__a21o_1 _09691_ (.A1(_02629_),
    .A2(_02630_),
    .B1(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__nand3_1 _09692_ (.A(_02629_),
    .B(_02630_),
    .C(_02631_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21bo_1 _09693_ (.A1(_01920_),
    .A2(_01922_),
    .B1_N(_01921_),
    .X(_02634_));
 sky130_fd_sc_hd__nand3_1 _09694_ (.A(_02632_),
    .B(_02633_),
    .C(_02634_),
    .Y(_02636_));
 sky130_fd_sc_hd__a21o_1 _09695_ (.A1(_02632_),
    .A2(_02633_),
    .B1(_02634_),
    .X(_02637_));
 sky130_fd_sc_hd__nand3_1 _09696_ (.A(_02628_),
    .B(_02636_),
    .C(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__a21o_1 _09697_ (.A1(_02636_),
    .A2(_02637_),
    .B1(_02628_),
    .X(_02639_));
 sky130_fd_sc_hd__a21bo_1 _09698_ (.A1(_01917_),
    .A2(_01926_),
    .B1_N(_01925_),
    .X(_02640_));
 sky130_fd_sc_hd__and3_1 _09699_ (.A(_02638_),
    .B(_02639_),
    .C(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__a21oi_1 _09700_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02640_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor3_1 _09701_ (.A(_02621_),
    .B(_02641_),
    .C(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__o21a_1 _09702_ (.A1(_02641_),
    .A2(_02642_),
    .B1(_02621_),
    .X(_02644_));
 sky130_fd_sc_hd__a211o_1 _09703_ (.A1(_02611_),
    .A2(_01932_),
    .B1(_02643_),
    .C1(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__o211ai_1 _09704_ (.A1(_02643_),
    .A2(_02644_),
    .B1(_02611_),
    .C1(_01932_),
    .Y(_02647_));
 sky130_fd_sc_hd__or4bb_2 _09705_ (.A(_02609_),
    .B(_02610_),
    .C_N(_02645_),
    .D_N(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__a2bb2o_1 _09706_ (.A1_N(_02609_),
    .A2_N(_02610_),
    .B1(_02645_),
    .B2(_02647_),
    .X(_02649_));
 sky130_fd_sc_hd__o211a_1 _09707_ (.A1(_02000_),
    .A2(_02585_),
    .B1(_02648_),
    .C1(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__a211oi_2 _09708_ (.A1(_02648_),
    .A2(_02649_),
    .B1(_02000_),
    .C1(_02585_),
    .Y(_02651_));
 sky130_fd_sc_hd__nor3_2 _09709_ (.A(_02584_),
    .B(_02650_),
    .C(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__o21a_1 _09710_ (.A1(_02650_),
    .A2(_02651_),
    .B1(_02584_),
    .X(_02653_));
 sky130_fd_sc_hd__a211o_1 _09711_ (.A1(_02582_),
    .A2(_02583_),
    .B1(_02652_),
    .C1(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__o211ai_4 _09712_ (.A1(_02652_),
    .A2(_02653_),
    .B1(_02582_),
    .C1(_02583_),
    .Y(_02655_));
 sky130_fd_sc_hd__nand3_2 _09713_ (.A(_02581_),
    .B(_02654_),
    .C(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21o_1 _09714_ (.A1(_02654_),
    .A2(_02655_),
    .B1(_02581_),
    .X(_02658_));
 sky130_fd_sc_hd__o211ai_4 _09715_ (.A1(_01961_),
    .A2(net293),
    .B1(_02656_),
    .C1(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__a211o_1 _09716_ (.A1(_02656_),
    .A2(_02658_),
    .B1(_01961_),
    .C1(_02579_),
    .X(_02660_));
 sky130_fd_sc_hd__nand3_2 _09717_ (.A(_02578_),
    .B(_02659_),
    .C(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__a21o_1 _09718_ (.A1(_02659_),
    .A2(_02660_),
    .B1(_02578_),
    .X(_02662_));
 sky130_fd_sc_hd__o211a_1 _09719_ (.A1(_02105_),
    .A2(_02107_),
    .B1(_02661_),
    .C1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__a211o_1 _09720_ (.A1(_02661_),
    .A2(_02662_),
    .B1(_02105_),
    .C1(_02107_),
    .X(_02664_));
 sky130_fd_sc_hd__and2b_1 _09721_ (.A_N(_02663_),
    .B(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__xor2_4 _09722_ (.A(_02453_),
    .B(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__a21bo_2 _09723_ (.A1(_02055_),
    .A2(_02102_),
    .B1_N(_02101_),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_2 _09724_ (.A(_02192_),
    .B(_02194_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_2 _09725_ (.A(_01996_),
    .B(_01999_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_01992_),
    .B(_01995_),
    .Y(_02671_));
 sky130_fd_sc_hd__o21bai_2 _09727_ (.A1(_02008_),
    .A2(_02016_),
    .B1_N(_02015_),
    .Y(_02672_));
 sky130_fd_sc_hd__or2_1 _09728_ (.A(_01989_),
    .B(_01991_),
    .X(_02673_));
 sky130_fd_sc_hd__a32oi_4 _09729_ (.A1(_05980_),
    .A2(net249),
    .A3(_02005_),
    .B1(_02004_),
    .B2(_00834_),
    .Y(_02674_));
 sky130_fd_sc_hd__a22oi_1 _09730_ (.A1(_05980_),
    .A2(_01367_),
    .B1(_01987_),
    .B2(_03853_),
    .Y(_02675_));
 sky130_fd_sc_hd__and4_2 _09731_ (.A(net236),
    .B(net237),
    .C(net250),
    .D(net251),
    .X(_02676_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(_02675_),
    .B(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__xor2_1 _09733_ (.A(_02674_),
    .B(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__xnor2_1 _09734_ (.A(_02673_),
    .B(_02678_),
    .Y(_02680_));
 sky130_fd_sc_hd__xnor2_1 _09735_ (.A(_02672_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor2_1 _09736_ (.A(_02671_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__a22o_1 _09737_ (.A1(_02030_),
    .A2(_02028_),
    .B1(_02032_),
    .B2(_02018_),
    .X(_02683_));
 sky130_fd_sc_hd__and2b_1 _09738_ (.A_N(_02682_),
    .B(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__or2b_1 _09739_ (.A(_02683_),
    .B_N(_02682_),
    .X(_02685_));
 sky130_fd_sc_hd__or2b_2 _09740_ (.A(_02684_),
    .B_N(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__xor2_4 _09741_ (.A(_02670_),
    .B(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__and3_1 _09742_ (.A(net247),
    .B(net239),
    .C(net248),
    .X(_02688_));
 sky130_fd_sc_hd__a22o_1 _09743_ (.A1(net239),
    .A2(net248),
    .B1(net240),
    .B2(net247),
    .X(_02689_));
 sky130_fd_sc_hd__a21bo_1 _09744_ (.A1(_01385_),
    .A2(_02688_),
    .B1_N(_02689_),
    .X(_02691_));
 sky130_fd_sc_hd__nand2_2 _09745_ (.A(_06384_),
    .B(_00830_),
    .Y(_02692_));
 sky130_fd_sc_hd__xor2_4 _09746_ (.A(_02691_),
    .B(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__buf_2 _09747_ (.A(net241),
    .X(_02694_));
 sky130_fd_sc_hd__buf_2 _09748_ (.A(net242),
    .X(_02695_));
 sky130_fd_sc_hd__a22oi_1 _09749_ (.A1(_05969_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_03864_),
    .Y(_02696_));
 sky130_fd_sc_hd__and4_1 _09750_ (.A(_03864_),
    .B(net246),
    .C(net241),
    .D(net242),
    .X(_02697_));
 sky130_fd_sc_hd__nor2_1 _09751_ (.A(_02696_),
    .B(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__a21bo_1 _09752_ (.A1(_02009_),
    .A2(_02011_),
    .B1_N(_02010_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_1 _09753_ (.A(_02698_),
    .B(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__or2_1 _09754_ (.A(_02698_),
    .B(_02699_),
    .X(_02702_));
 sky130_fd_sc_hd__and2b_1 _09755_ (.A_N(_02700_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__xor2_2 _09756_ (.A(_02693_),
    .B(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__nand2_1 _09757_ (.A(_02021_),
    .B(_02023_),
    .Y(_02705_));
 sky130_fd_sc_hd__a21bo_1 _09758_ (.A1(_02036_),
    .A2(_02039_),
    .B1_N(_02037_),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _09759_ (.A1(_06375_),
    .A2(net11),
    .B1(net13),
    .B2(net254),
    .X(_02707_));
 sky130_fd_sc_hd__nand4_2 _09760_ (.A(net254),
    .B(_06375_),
    .C(net11),
    .D(net13),
    .Y(_02708_));
 sky130_fd_sc_hd__a22o_1 _09761_ (.A1(_03820_),
    .A2(net14),
    .B1(_02707_),
    .B2(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__nand4_2 _09762_ (.A(_03820_),
    .B(_02019_),
    .C(_02707_),
    .D(_02708_),
    .Y(_02710_));
 sky130_fd_sc_hd__nand3_1 _09763_ (.A(_02706_),
    .B(_02709_),
    .C(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a21o_1 _09764_ (.A1(_02709_),
    .A2(_02710_),
    .B1(_02706_),
    .X(_02713_));
 sky130_fd_sc_hd__nand3_1 _09765_ (.A(_02705_),
    .B(_02711_),
    .C(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__a21o_1 _09766_ (.A1(_02711_),
    .A2(_02713_),
    .B1(_02705_),
    .X(_02715_));
 sky130_fd_sc_hd__a211o_1 _09767_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_02024_),
    .C1(_02025_),
    .X(_02716_));
 sky130_fd_sc_hd__o21a_1 _09768_ (.A1(_02029_),
    .A2(_02027_),
    .B1(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__nand3_1 _09769_ (.A(_02714_),
    .B(_02715_),
    .C(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21o_1 _09770_ (.A1(_02714_),
    .A2(_02715_),
    .B1(_02717_),
    .X(_02719_));
 sky130_fd_sc_hd__and3_1 _09771_ (.A(_02704_),
    .B(_02718_),
    .C(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__a21oi_1 _09772_ (.A1(_02718_),
    .A2(_02719_),
    .B1(_02704_),
    .Y(_02721_));
 sky130_fd_sc_hd__nor2_2 _09773_ (.A(_02720_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__a2bb2o_2 _09774_ (.A1_N(_02046_),
    .A2_N(_02040_),
    .B1(_01412_),
    .B2(_02043_),
    .X(_02724_));
 sky130_fd_sc_hd__a21oi_2 _09775_ (.A1(_02081_),
    .A2(_02088_),
    .B1(_02087_),
    .Y(_02725_));
 sky130_fd_sc_hd__a22o_1 _09776_ (.A1(net9),
    .A2(net3),
    .B1(net4),
    .B2(_05882_),
    .X(_02726_));
 sky130_fd_sc_hd__nand4_4 _09777_ (.A(_05882_),
    .B(_06368_),
    .C(_00850_),
    .D(net4),
    .Y(_02727_));
 sky130_fd_sc_hd__a22o_1 _09778_ (.A1(_00357_),
    .A2(_00822_),
    .B1(_02726_),
    .B2(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__nand4_4 _09779_ (.A(_00357_),
    .B(_00822_),
    .C(_02726_),
    .D(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _09780_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__clkbuf_4 _09781_ (.A(net5),
    .X(_02731_));
 sky130_fd_sc_hd__a22oi_2 _09782_ (.A1(_03732_),
    .A2(net66),
    .B1(_02731_),
    .B2(_03798_),
    .Y(_02732_));
 sky130_fd_sc_hd__and4_2 _09783_ (.A(net51),
    .B(_03798_),
    .C(net66),
    .D(net5),
    .X(_02733_));
 sky130_fd_sc_hd__nor2_1 _09784_ (.A(_02732_),
    .B(_02733_),
    .Y(_02735_));
 sky130_fd_sc_hd__o21bai_2 _09785_ (.A1(_02042_),
    .A2(_02044_),
    .B1_N(_02041_),
    .Y(_02736_));
 sky130_fd_sc_hd__xnor2_2 _09786_ (.A(_02735_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__xnor2_2 _09787_ (.A(_02730_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__xnor2_2 _09788_ (.A(_02725_),
    .B(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__xor2_4 _09789_ (.A(_02724_),
    .B(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__nor2_1 _09790_ (.A(_02035_),
    .B(_02047_),
    .Y(_02741_));
 sky130_fd_sc_hd__a21oi_4 _09791_ (.A1(_02034_),
    .A2(_02048_),
    .B1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__xnor2_4 _09792_ (.A(_02740_),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__xnor2_4 _09793_ (.A(_02722_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__and2b_1 _09794_ (.A_N(_02050_),
    .B(_02049_),
    .X(_02746_));
 sky130_fd_sc_hd__a21oi_2 _09795_ (.A1(_02033_),
    .A2(_02051_),
    .B1(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_4 _09796_ (.A(_02744_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__xor2_4 _09797_ (.A(_02687_),
    .B(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__or2_1 _09798_ (.A(_02093_),
    .B(_02095_),
    .X(_02750_));
 sky130_fd_sc_hd__a21boi_2 _09799_ (.A1(_02126_),
    .A2(_02156_),
    .B1_N(_02155_),
    .Y(_02751_));
 sky130_fd_sc_hd__or2_2 _09800_ (.A(_02079_),
    .B(_02091_),
    .X(_02752_));
 sky130_fd_sc_hd__a21oi_2 _09801_ (.A1(_02113_),
    .A2(_02124_),
    .B1(_02123_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _09802_ (.A(_02084_),
    .B(_02086_),
    .Y(_02754_));
 sky130_fd_sc_hd__a32o_1 _09803_ (.A1(_06347_),
    .A2(_00387_),
    .A3(_02073_),
    .B1(_02072_),
    .B2(_01444_),
    .X(_02755_));
 sky130_fd_sc_hd__a22o_1 _09804_ (.A1(net54),
    .A2(net63),
    .B1(net64),
    .B2(net53),
    .X(_02757_));
 sky130_fd_sc_hd__nand4_2 _09805_ (.A(net53),
    .B(net54),
    .C(_00397_),
    .D(_00872_),
    .Y(_02758_));
 sky130_fd_sc_hd__a22o_1 _09806_ (.A1(_05750_),
    .A2(net65),
    .B1(_02757_),
    .B2(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__nand4_2 _09807_ (.A(_05750_),
    .B(_01434_),
    .C(_02757_),
    .D(_02758_),
    .Y(_02760_));
 sky130_fd_sc_hd__and3_1 _09808_ (.A(_02755_),
    .B(_02759_),
    .C(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__a21o_1 _09809_ (.A1(_02759_),
    .A2(_02760_),
    .B1(_02755_),
    .X(_02762_));
 sky130_fd_sc_hd__and2b_1 _09810_ (.A_N(_02761_),
    .B(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__xnor2_2 _09811_ (.A(_02754_),
    .B(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__clkbuf_4 _09812_ (.A(net58),
    .X(_02765_));
 sky130_fd_sc_hd__and3_1 _09813_ (.A(net60),
    .B(net61),
    .C(net57),
    .X(_02766_));
 sky130_fd_sc_hd__a22o_1 _09814_ (.A1(net61),
    .A2(net57),
    .B1(net58),
    .B2(net60),
    .X(_02768_));
 sky130_fd_sc_hd__a21bo_1 _09815_ (.A1(_02765_),
    .A2(_02766_),
    .B1_N(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__nand2_1 _09816_ (.A(_06347_),
    .B(_00879_),
    .Y(_02770_));
 sky130_fd_sc_hd__xnor2_2 _09817_ (.A(_02769_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__a22oi_1 _09818_ (.A1(_05498_),
    .A2(_01443_),
    .B1(_02064_),
    .B2(_03579_),
    .Y(_02772_));
 sky130_fd_sc_hd__and4_1 _09819_ (.A(net69),
    .B(_05498_),
    .C(net83),
    .D(net84),
    .X(_02773_));
 sky130_fd_sc_hd__nor2_1 _09820_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__a21bo_1 _09821_ (.A1(_02065_),
    .A2(_02067_),
    .B1_N(_02066_),
    .X(_02775_));
 sky130_fd_sc_hd__xor2_1 _09822_ (.A(_02774_),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__xnor2_2 _09823_ (.A(_02771_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__a21boi_2 _09824_ (.A1(_02071_),
    .A2(_02076_),
    .B1_N(_02070_),
    .Y(_02779_));
 sky130_fd_sc_hd__xnor2_2 _09825_ (.A(_02777_),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__xnor2_2 _09826_ (.A(_02764_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__xnor2_2 _09827_ (.A(_02753_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__xnor2_2 _09828_ (.A(_02752_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__xor2_2 _09829_ (.A(_02751_),
    .B(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__xnor2_1 _09830_ (.A(_02750_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__a21boi_1 _09831_ (.A1(_02059_),
    .A2(_02098_),
    .B1_N(_02097_),
    .Y(_02786_));
 sky130_fd_sc_hd__nor2_1 _09832_ (.A(_02785_),
    .B(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_1 _09833_ (.A(_02785_),
    .B(_02786_),
    .Y(_02788_));
 sky130_fd_sc_hd__and2b_1 _09834_ (.A_N(_02787_),
    .B(_02788_),
    .X(_02790_));
 sky130_fd_sc_hd__xnor2_4 _09835_ (.A(_02749_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__xnor2_4 _09836_ (.A(_02669_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__xor2_4 _09837_ (.A(_02667_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__inv_2 _09838_ (.A(_02188_),
    .Y(_02794_));
 sky130_fd_sc_hd__or2_2 _09839_ (.A(_02794_),
    .B(_02190_),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(_02119_),
    .B(_02121_),
    .Y(_02796_));
 sky130_fd_sc_hd__a21bo_1 _09841_ (.A1(_02131_),
    .A2(_02138_),
    .B1_N(_02137_),
    .X(_02797_));
 sky130_fd_sc_hd__a41o_1 _09842_ (.A1(_06424_),
    .A2(_06410_),
    .A3(_00431_),
    .A4(_00421_),
    .B1(_02118_),
    .X(_02798_));
 sky130_fd_sc_hd__buf_2 _09843_ (.A(net75),
    .X(_02799_));
 sky130_fd_sc_hd__a32o_1 _09844_ (.A1(net79),
    .A2(_01487_),
    .A3(_02128_),
    .B1(_02127_),
    .B2(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__a22o_1 _09845_ (.A1(net72),
    .A2(_00421_),
    .B1(net73),
    .B2(_06410_),
    .X(_02802_));
 sky130_fd_sc_hd__nand4_1 _09846_ (.A(_06410_),
    .B(_00431_),
    .C(_00421_),
    .D(_01487_),
    .Y(_02803_));
 sky130_fd_sc_hd__a22o_1 _09847_ (.A1(_06424_),
    .A2(_00937_),
    .B1(_02802_),
    .B2(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__nand4_1 _09848_ (.A(_06424_),
    .B(_00937_),
    .C(_02802_),
    .D(_02803_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand3_1 _09849_ (.A(_02801_),
    .B(_02804_),
    .C(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__a21o_1 _09850_ (.A1(_02804_),
    .A2(_02805_),
    .B1(_02801_),
    .X(_02807_));
 sky130_fd_sc_hd__nand3_1 _09851_ (.A(_02798_),
    .B(_02806_),
    .C(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__a21o_1 _09852_ (.A1(_02806_),
    .A2(_02807_),
    .B1(_02798_),
    .X(_02809_));
 sky130_fd_sc_hd__and3_1 _09853_ (.A(_02797_),
    .B(_02808_),
    .C(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a21o_1 _09854_ (.A1(_02808_),
    .A2(_02809_),
    .B1(_02797_),
    .X(_02812_));
 sky130_fd_sc_hd__or2b_1 _09855_ (.A(_02810_),
    .B_N(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__xnor2_2 _09856_ (.A(_02796_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__and3_1 _09857_ (.A(_02148_),
    .B(_02149_),
    .C(_02150_),
    .X(_02815_));
 sky130_fd_sc_hd__a22oi_1 _09858_ (.A1(net79),
    .A2(_01488_),
    .B1(_02799_),
    .B2(_03590_),
    .Y(_02816_));
 sky130_fd_sc_hd__and4_1 _09859_ (.A(_03590_),
    .B(net79),
    .C(_01488_),
    .D(net75),
    .X(_02817_));
 sky130_fd_sc_hd__nor2_1 _09860_ (.A(_02816_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__and4_1 _09861_ (.A(net104),
    .B(net105),
    .C(_00910_),
    .D(net119),
    .X(_02819_));
 sky130_fd_sc_hd__and4_1 _09862_ (.A(net103),
    .B(net120),
    .C(_02133_),
    .D(_02134_),
    .X(_02820_));
 sky130_fd_sc_hd__a22o_1 _09863_ (.A1(net106),
    .A2(net118),
    .B1(net119),
    .B2(net105),
    .X(_02821_));
 sky130_fd_sc_hd__nand4_2 _09864_ (.A(net105),
    .B(net106),
    .C(net118),
    .D(net119),
    .Y(_02823_));
 sky130_fd_sc_hd__a22o_1 _09865_ (.A1(net104),
    .A2(net120),
    .B1(_02821_),
    .B2(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__nand4_2 _09866_ (.A(net104),
    .B(_02132_),
    .C(_02821_),
    .D(_02823_),
    .Y(_02825_));
 sky130_fd_sc_hd__o211a_1 _09867_ (.A1(_02819_),
    .A2(_02820_),
    .B1(_02824_),
    .C1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__a211o_1 _09868_ (.A1(_02824_),
    .A2(_02825_),
    .B1(_02819_),
    .C1(_02820_),
    .X(_02827_));
 sky130_fd_sc_hd__and2b_1 _09869_ (.A_N(_02826_),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__xnor2_1 _09870_ (.A(_02818_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _09871_ (.A(_02143_),
    .B(_02145_),
    .Y(_02830_));
 sky130_fd_sc_hd__a32o_1 _09872_ (.A1(net114),
    .A2(net109),
    .A3(_02166_),
    .B1(_02165_),
    .B2(net110),
    .X(_02831_));
 sky130_fd_sc_hd__a22o_1 _09873_ (.A1(net116),
    .A2(net108),
    .B1(net109),
    .B2(net115),
    .X(_02832_));
 sky130_fd_sc_hd__nand4_1 _09874_ (.A(net115),
    .B(net116),
    .C(net108),
    .D(net109),
    .Y(_02834_));
 sky130_fd_sc_hd__and2_1 _09875_ (.A(net107),
    .B(net117),
    .X(_02835_));
 sky130_fd_sc_hd__a21o_1 _09876_ (.A1(_02832_),
    .A2(_02834_),
    .B1(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__nand3_1 _09877_ (.A(_02832_),
    .B(_02834_),
    .C(_02835_),
    .Y(_02837_));
 sky130_fd_sc_hd__nand3_1 _09878_ (.A(_02831_),
    .B(_02836_),
    .C(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21o_1 _09879_ (.A1(_02836_),
    .A2(_02837_),
    .B1(_02831_),
    .X(_02839_));
 sky130_fd_sc_hd__nand3_1 _09880_ (.A(_02830_),
    .B(_02838_),
    .C(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__a21o_1 _09881_ (.A1(_02838_),
    .A2(_02839_),
    .B1(_02830_),
    .X(_02841_));
 sky130_fd_sc_hd__a21bo_1 _09882_ (.A1(_02141_),
    .A2(_02147_),
    .B1_N(_02146_),
    .X(_02842_));
 sky130_fd_sc_hd__and3_1 _09883_ (.A(_02840_),
    .B(_02841_),
    .C(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a21oi_1 _09884_ (.A1(_02840_),
    .A2(_02841_),
    .B1(_02842_),
    .Y(_02845_));
 sky130_fd_sc_hd__or3_2 _09885_ (.A(_02829_),
    .B(_02843_),
    .C(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__o21ai_1 _09886_ (.A1(_02843_),
    .A2(_02845_),
    .B1(_02829_),
    .Y(_02847_));
 sky130_fd_sc_hd__o211a_1 _09887_ (.A1(_02815_),
    .A2(_02153_),
    .B1(_02846_),
    .C1(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__inv_2 _09888_ (.A(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__a211o_1 _09889_ (.A1(_02846_),
    .A2(_02847_),
    .B1(_02815_),
    .C1(_02153_),
    .X(_02850_));
 sky130_fd_sc_hd__and3_1 _09890_ (.A(_02814_),
    .B(_02849_),
    .C(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__a21oi_2 _09891_ (.A1(_02849_),
    .A2(_02850_),
    .B1(_02814_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand3_1 _09892_ (.A(_02159_),
    .B(_02183_),
    .C(_02184_),
    .Y(_02853_));
 sky130_fd_sc_hd__a31o_1 _09893_ (.A1(_01559_),
    .A2(_02177_),
    .A3(_02178_),
    .B1(_02181_),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _09894_ (.A(_02175_),
    .B(_02177_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21o_1 _09895_ (.A1(_02202_),
    .A2(_02209_),
    .B1(_02208_),
    .X(_02857_));
 sky130_fd_sc_hd__a22oi_1 _09896_ (.A1(_03381_),
    .A2(net181),
    .B1(_02164_),
    .B2(_03546_),
    .Y(_02858_));
 sky130_fd_sc_hd__and4_2 _09897_ (.A(net89),
    .B(net114),
    .C(net181),
    .D(net110),
    .X(_02859_));
 sky130_fd_sc_hd__nor2_2 _09898_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__and4_1 _09899_ (.A(net100),
    .B(_00059_),
    .C(_00453_),
    .D(_00953_),
    .X(_02861_));
 sky130_fd_sc_hd__and4_1 _09900_ (.A(net89),
    .B(_01524_),
    .C(_02170_),
    .D(_02171_),
    .X(_02862_));
 sky130_fd_sc_hd__a22o_1 _09901_ (.A1(net123),
    .A2(net177),
    .B1(net178),
    .B2(net111),
    .X(_02863_));
 sky130_fd_sc_hd__nand4_2 _09902_ (.A(net111),
    .B(net123),
    .C(net177),
    .D(net178),
    .Y(_02864_));
 sky130_fd_sc_hd__and2_1 _09903_ (.A(net100),
    .B(net180),
    .X(_02865_));
 sky130_fd_sc_hd__a21o_1 _09904_ (.A1(_02863_),
    .A2(_02864_),
    .B1(_02865_),
    .X(_02867_));
 sky130_fd_sc_hd__nand3_1 _09905_ (.A(_02863_),
    .B(_02864_),
    .C(_02865_),
    .Y(_02868_));
 sky130_fd_sc_hd__o211ai_2 _09906_ (.A1(_02861_),
    .A2(_02862_),
    .B1(_02867_),
    .C1(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__a211o_1 _09907_ (.A1(_02867_),
    .A2(_02868_),
    .B1(_02861_),
    .C1(_02862_),
    .X(_02870_));
 sky130_fd_sc_hd__nand3_2 _09908_ (.A(_02860_),
    .B(_02869_),
    .C(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__a21o_1 _09909_ (.A1(_02869_),
    .A2(_02870_),
    .B1(_02860_),
    .X(_02872_));
 sky130_fd_sc_hd__nand3_4 _09910_ (.A(_02857_),
    .B(_02871_),
    .C(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__a21o_1 _09911_ (.A1(_02871_),
    .A2(_02872_),
    .B1(_02857_),
    .X(_02874_));
 sky130_fd_sc_hd__nand3_4 _09912_ (.A(_02856_),
    .B(_02873_),
    .C(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__a21o_1 _09913_ (.A1(_02873_),
    .A2(_02874_),
    .B1(_02856_),
    .X(_02876_));
 sky130_fd_sc_hd__o211ai_4 _09914_ (.A1(_02231_),
    .A2(net304),
    .B1(_02875_),
    .C1(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__a211o_1 _09915_ (.A1(_02875_),
    .A2(_02876_),
    .B1(_02231_),
    .C1(net304),
    .X(_02879_));
 sky130_fd_sc_hd__and3_1 _09916_ (.A(_02854_),
    .B(_02878_),
    .C(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__a21oi_1 _09917_ (.A1(_02878_),
    .A2(_02879_),
    .B1(_02854_),
    .Y(_02881_));
 sky130_fd_sc_hd__a211o_1 _09918_ (.A1(_02183_),
    .A2(_02853_),
    .B1(_02880_),
    .C1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__o211ai_1 _09919_ (.A1(_02880_),
    .A2(_02881_),
    .B1(_02183_),
    .C1(_02853_),
    .Y(_02883_));
 sky130_fd_sc_hd__or4bb_2 _09920_ (.A(_02851_),
    .B(_02852_),
    .C_N(_02882_),
    .D_N(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__a2bb2o_1 _09921_ (.A1_N(_02851_),
    .A2_N(_02852_),
    .B1(_02882_),
    .B2(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__o211a_1 _09922_ (.A1(_02259_),
    .A2(_02261_),
    .B1(_02884_),
    .C1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__a211o_1 _09923_ (.A1(_02884_),
    .A2(_02885_),
    .B1(_02259_),
    .C1(_02261_),
    .X(_02887_));
 sky130_fd_sc_hd__or2b_2 _09924_ (.A(_02886_),
    .B_N(_02887_),
    .X(_02889_));
 sky130_fd_sc_hd__xnor2_4 _09925_ (.A(_02795_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__a21bo_1 _09926_ (.A1(_02266_),
    .A2(_02299_),
    .B1_N(_02298_),
    .X(_02891_));
 sky130_fd_sc_hd__nand2_1 _09927_ (.A(_02204_),
    .B(_02206_),
    .Y(_02892_));
 sky130_fd_sc_hd__o21bai_1 _09928_ (.A1(_02212_),
    .A2(_02216_),
    .B1_N(_02213_),
    .Y(_02893_));
 sky130_fd_sc_hd__a22oi_1 _09929_ (.A1(net175),
    .A2(net145),
    .B1(net156),
    .B2(net174),
    .Y(_02894_));
 sky130_fd_sc_hd__and4_1 _09930_ (.A(net174),
    .B(net175),
    .C(net145),
    .D(net156),
    .X(_02895_));
 sky130_fd_sc_hd__a2bb2o_1 _09931_ (.A1_N(_02894_),
    .A2_N(_02895_),
    .B1(net176),
    .B2(_00985_),
    .X(_02896_));
 sky130_fd_sc_hd__or4bb_1 _09932_ (.A(_02894_),
    .B(_02895_),
    .C_N(net176),
    .D_N(_00985_),
    .X(_02897_));
 sky130_fd_sc_hd__nand3_1 _09933_ (.A(_02893_),
    .B(_02896_),
    .C(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__a21o_1 _09934_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_02893_),
    .X(_02900_));
 sky130_fd_sc_hd__and3_1 _09935_ (.A(_02892_),
    .B(_02898_),
    .C(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__a21oi_1 _09936_ (.A1(_02898_),
    .A2(_02900_),
    .B1(_02892_),
    .Y(_02902_));
 sky130_fd_sc_hd__nor2_1 _09937_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__buf_2 _09938_ (.A(net198),
    .X(_02904_));
 sky130_fd_sc_hd__a22oi_1 _09939_ (.A1(_05115_),
    .A2(_01562_),
    .B1(_02904_),
    .B2(_03337_),
    .Y(_02905_));
 sky130_fd_sc_hd__and4_2 _09940_ (.A(net183),
    .B(net184),
    .C(net197),
    .D(net198),
    .X(_02906_));
 sky130_fd_sc_hd__nor2_1 _09941_ (.A(_02905_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__and4_1 _09942_ (.A(_00047_),
    .B(_00058_),
    .C(_00489_),
    .D(_00481_),
    .X(_02908_));
 sky130_fd_sc_hd__and4_1 _09943_ (.A(net184),
    .B(net196),
    .C(_02221_),
    .D(_02222_),
    .X(_02909_));
 sky130_fd_sc_hd__a22o_1 _09944_ (.A1(net186),
    .A2(net195),
    .B1(net187),
    .B2(_00989_),
    .X(_02911_));
 sky130_fd_sc_hd__nand4_1 _09945_ (.A(_00989_),
    .B(net186),
    .C(_00480_),
    .D(net187),
    .Y(_02912_));
 sky130_fd_sc_hd__a22o_1 _09946_ (.A1(_00047_),
    .A2(_01567_),
    .B1(_02911_),
    .B2(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__nand4_1 _09947_ (.A(_00049_),
    .B(_01567_),
    .C(_02911_),
    .D(_02912_),
    .Y(_02914_));
 sky130_fd_sc_hd__o211ai_2 _09948_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_02913_),
    .C1(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__a211o_1 _09949_ (.A1(_02913_),
    .A2(_02914_),
    .B1(_02908_),
    .C1(_02909_),
    .X(_02916_));
 sky130_fd_sc_hd__nand3_2 _09950_ (.A(_02907_),
    .B(_02915_),
    .C(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21o_1 _09951_ (.A1(_02915_),
    .A2(_02916_),
    .B1(_02907_),
    .X(_02918_));
 sky130_fd_sc_hd__a21bo_1 _09952_ (.A1(_02217_),
    .A2(_02226_),
    .B1_N(_02225_),
    .X(_02919_));
 sky130_fd_sc_hd__nand3_4 _09953_ (.A(_02917_),
    .B(_02918_),
    .C(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__a21o_1 _09954_ (.A1(_02917_),
    .A2(_02918_),
    .B1(_02919_),
    .X(_02922_));
 sky130_fd_sc_hd__nand3_2 _09955_ (.A(_02903_),
    .B(_02920_),
    .C(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21o_1 _09956_ (.A1(_02920_),
    .A2(_02922_),
    .B1(_02903_),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_2 _09957_ (.A(_02923_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_2 _09958_ (.A(_02244_),
    .B(_02246_),
    .Y(_02926_));
 sky130_fd_sc_hd__o211a_1 _09959_ (.A1(_02276_),
    .A2(_02277_),
    .B1(_01610_),
    .C1(_01611_),
    .X(_02927_));
 sky130_fd_sc_hd__a211o_1 _09960_ (.A1(_01610_),
    .A2(_01611_),
    .B1(_02276_),
    .C1(_02277_),
    .X(_02928_));
 sky130_fd_sc_hd__o21a_1 _09961_ (.A1(_02272_),
    .A2(_02927_),
    .B1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_02241_),
    .B(_02243_),
    .Y(_02930_));
 sky130_fd_sc_hd__o21bai_2 _09963_ (.A1(_02268_),
    .A2(_02271_),
    .B1_N(_02269_),
    .Y(_02931_));
 sky130_fd_sc_hd__nand2_1 _09964_ (.A(net192),
    .B(net189),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _09965_ (.A(net193),
    .B(net188),
    .Y(_02934_));
 sky130_fd_sc_hd__xor2_2 _09966_ (.A(_02933_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__xor2_2 _09967_ (.A(_02931_),
    .B(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__xnor2_2 _09968_ (.A(_02930_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__xor2_2 _09969_ (.A(_02929_),
    .B(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__xor2_2 _09970_ (.A(_02926_),
    .B(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__a21boi_2 _09971_ (.A1(_02235_),
    .A2(_02249_),
    .B1_N(_02248_),
    .Y(_02940_));
 sky130_fd_sc_hd__xor2_2 _09972_ (.A(_02939_),
    .B(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__xor2_1 _09973_ (.A(_02925_),
    .B(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__xnor2_1 _09974_ (.A(_02891_),
    .B(_02942_),
    .Y(_02944_));
 sky130_fd_sc_hd__a21oi_2 _09975_ (.A1(_02255_),
    .A2(_02257_),
    .B1(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__and3_1 _09976_ (.A(_02255_),
    .B(_02257_),
    .C(_02944_),
    .X(_02946_));
 sky130_fd_sc_hd__nor2_2 _09977_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__a31o_2 _09978_ (.A1(_02290_),
    .A2(_02291_),
    .A3(_02292_),
    .B1(_02296_),
    .X(_02948_));
 sky130_fd_sc_hd__o21bai_2 _09979_ (.A1(_02303_),
    .A2(_02323_),
    .B1_N(_02322_),
    .Y(_02949_));
 sky130_fd_sc_hd__and3_1 _09980_ (.A(net219),
    .B(net220),
    .C(net232),
    .X(_02950_));
 sky130_fd_sc_hd__a22oi_1 _09981_ (.A1(net220),
    .A2(net231),
    .B1(net232),
    .B2(net219),
    .Y(_02951_));
 sky130_fd_sc_hd__a21oi_2 _09982_ (.A1(_01023_),
    .A2(_02950_),
    .B1(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__and2_1 _09983_ (.A(net218),
    .B(net233),
    .X(_02953_));
 sky130_fd_sc_hd__xnor2_2 _09984_ (.A(_02952_),
    .B(_02953_),
    .Y(_02955_));
 sky130_fd_sc_hd__and4_1 _09985_ (.A(_04741_),
    .B(_00086_),
    .C(_00507_),
    .D(_01034_),
    .X(_02956_));
 sky130_fd_sc_hd__a22o_1 _09986_ (.A1(net229),
    .A2(net222),
    .B1(net224),
    .B2(net228),
    .X(_02957_));
 sky130_fd_sc_hd__nand4_1 _09987_ (.A(net228),
    .B(net229),
    .C(net222),
    .D(net224),
    .Y(_02958_));
 sky130_fd_sc_hd__and2_1 _09988_ (.A(net221),
    .B(net230),
    .X(_02959_));
 sky130_fd_sc_hd__a21o_1 _09989_ (.A1(_02957_),
    .A2(_02958_),
    .B1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__nand3_1 _09990_ (.A(_02957_),
    .B(_02958_),
    .C(_02959_),
    .Y(_02961_));
 sky130_fd_sc_hd__o211ai_2 _09991_ (.A1(_02956_),
    .A2(_02277_),
    .B1(_02960_),
    .C1(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__a211o_1 _09992_ (.A1(_02960_),
    .A2(_02961_),
    .B1(_02956_),
    .C1(_02277_),
    .X(_02963_));
 sky130_fd_sc_hd__nand2_1 _09993_ (.A(_02962_),
    .B(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__xor2_2 _09994_ (.A(_02955_),
    .B(_02964_),
    .X(_02966_));
 sky130_fd_sc_hd__nand2_1 _09995_ (.A(_02283_),
    .B(_02287_),
    .Y(_02967_));
 sky130_fd_sc_hd__o21bai_2 _09996_ (.A1(_02304_),
    .A2(_02308_),
    .B1_N(_02305_),
    .Y(_02968_));
 sky130_fd_sc_hd__and4_2 _09997_ (.A(net33),
    .B(net227),
    .C(net49),
    .D(net225),
    .X(_02969_));
 sky130_fd_sc_hd__a22o_1 _09998_ (.A1(_03084_),
    .A2(net49),
    .B1(net225),
    .B2(net227),
    .X(_02970_));
 sky130_fd_sc_hd__or2b_1 _09999_ (.A(_02969_),
    .B_N(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__xnor2_2 _10000_ (.A(_02968_),
    .B(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__xor2_2 _10001_ (.A(_02967_),
    .B(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__o21ba_1 _10002_ (.A1(_01619_),
    .A2(_02289_),
    .B1_N(_02288_),
    .X(_02974_));
 sky130_fd_sc_hd__xnor2_2 _10003_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__xnor2_2 _10004_ (.A(_02966_),
    .B(_02975_),
    .Y(_02977_));
 sky130_fd_sc_hd__xnor2_2 _10005_ (.A(_02949_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__xor2_4 _10006_ (.A(_02948_),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__nand2_2 _10007_ (.A(_02318_),
    .B(_02320_),
    .Y(_02980_));
 sky130_fd_sc_hd__a21o_1 _10008_ (.A1(_01655_),
    .A2(_02335_),
    .B1(_02334_),
    .X(_02981_));
 sky130_fd_sc_hd__a22oi_4 _10009_ (.A1(net37),
    .A2(net46),
    .B1(_01051_),
    .B2(net36),
    .Y(_02982_));
 sky130_fd_sc_hd__and4_1 _10010_ (.A(net36),
    .B(net37),
    .C(net46),
    .D(net47),
    .X(_02983_));
 sky130_fd_sc_hd__or2_1 _10011_ (.A(_02982_),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__nand2_2 _10012_ (.A(_04906_),
    .B(net48),
    .Y(_02985_));
 sky130_fd_sc_hd__xnor2_1 _10013_ (.A(_02984_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__a22o_1 _10014_ (.A1(net43),
    .A2(net39),
    .B1(net40),
    .B2(net42),
    .X(_02988_));
 sky130_fd_sc_hd__nand4_2 _10015_ (.A(_03194_),
    .B(_04862_),
    .C(net39),
    .D(net40),
    .Y(_02989_));
 sky130_fd_sc_hd__and2_1 _10016_ (.A(net44),
    .B(net38),
    .X(_02990_));
 sky130_fd_sc_hd__a21o_1 _10017_ (.A1(_02988_),
    .A2(_02989_),
    .B1(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__nand3_1 _10018_ (.A(_02988_),
    .B(_02989_),
    .C(_02990_),
    .Y(_02992_));
 sky130_fd_sc_hd__a21bo_1 _10019_ (.A1(_02312_),
    .A2(_02314_),
    .B1_N(_02313_),
    .X(_02993_));
 sky130_fd_sc_hd__and3_1 _10020_ (.A(_02991_),
    .B(_02992_),
    .C(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__a21oi_1 _10021_ (.A1(_02991_),
    .A2(_02992_),
    .B1(_02993_),
    .Y(_02995_));
 sky130_fd_sc_hd__or3_1 _10022_ (.A(_02986_),
    .B(_02994_),
    .C(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__o21ai_1 _10023_ (.A1(_02994_),
    .A2(_02995_),
    .B1(_02986_),
    .Y(_02997_));
 sky130_fd_sc_hd__and3_1 _10024_ (.A(_02981_),
    .B(_02996_),
    .C(_02997_),
    .X(_02999_));
 sky130_fd_sc_hd__a21o_1 _10025_ (.A1(_02996_),
    .A2(_02997_),
    .B1(_02981_),
    .X(_03000_));
 sky130_fd_sc_hd__or2b_2 _10026_ (.A(_02999_),
    .B_N(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__xnor2_4 _10027_ (.A(_02980_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand2_1 _10028_ (.A(_02331_),
    .B(_02333_),
    .Y(_03003_));
 sky130_fd_sc_hd__a31o_1 _10029_ (.A1(_04939_),
    .A2(net45),
    .A3(_02340_),
    .B1(_02338_),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_1 _10030_ (.A1(_04939_),
    .A2(net56),
    .B1(net67),
    .B2(_03095_),
    .X(_03005_));
 sky130_fd_sc_hd__buf_2 _10031_ (.A(net67),
    .X(_03006_));
 sky130_fd_sc_hd__nand4_1 _10032_ (.A(_03095_),
    .B(_04939_),
    .C(net56),
    .D(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_03005_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__xnor2_1 _10034_ (.A(_03004_),
    .B(_03008_),
    .Y(_03010_));
 sky130_fd_sc_hd__and2_1 _10035_ (.A(_03003_),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(_03003_),
    .B(_03010_),
    .Y(_03012_));
 sky130_fd_sc_hd__nor2_2 _10037_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__and3_1 _10038_ (.A(net23),
    .B(net201),
    .C(net34),
    .X(_03014_));
 sky130_fd_sc_hd__a22o_1 _10039_ (.A1(net201),
    .A2(net34),
    .B1(net212),
    .B2(net23),
    .X(_03015_));
 sky130_fd_sc_hd__a21bo_2 _10040_ (.A1(_01666_),
    .A2(_03014_),
    .B1_N(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__nand2_2 _10041_ (.A(_00549_),
    .B(_01072_),
    .Y(_03017_));
 sky130_fd_sc_hd__xor2_4 _10042_ (.A(_03016_),
    .B(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_4 _10043_ (.A(net234),
    .X(_03019_));
 sky130_fd_sc_hd__a22oi_1 _10044_ (.A1(net12),
    .A2(_01667_),
    .B1(_03019_),
    .B2(_03106_),
    .Y(_03021_));
 sky130_fd_sc_hd__and4_1 _10045_ (.A(_03106_),
    .B(net12),
    .C(net223),
    .D(net234),
    .X(_03022_));
 sky130_fd_sc_hd__nor2_2 _10046_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__a21bo_1 _10047_ (.A1(_02344_),
    .A2(_02346_),
    .B1_N(_02345_),
    .X(_03024_));
 sky130_fd_sc_hd__xor2_4 _10048_ (.A(_03023_),
    .B(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__xor2_4 _10049_ (.A(_03018_),
    .B(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__a21bo_2 _10050_ (.A1(_02343_),
    .A2(_02352_),
    .B1_N(_02351_),
    .X(_03027_));
 sky130_fd_sc_hd__xor2_4 _10051_ (.A(_03026_),
    .B(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__xor2_4 _10052_ (.A(_03013_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o21bai_4 _10053_ (.A1(_02337_),
    .A2(_02357_),
    .B1_N(_02356_),
    .Y(_03030_));
 sky130_fd_sc_hd__xor2_4 _10054_ (.A(_03029_),
    .B(_03030_),
    .X(_03032_));
 sky130_fd_sc_hd__xor2_4 _10055_ (.A(_03002_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__o211a_1 _10056_ (.A1(_02326_),
    .A2(_01680_),
    .B1(_02358_),
    .C1(_02359_),
    .X(_03034_));
 sky130_fd_sc_hd__a21oi_4 _10057_ (.A1(_02325_),
    .A2(_02362_),
    .B1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_4 _10058_ (.A(_03033_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__xor2_4 _10059_ (.A(_02979_),
    .B(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__a211oi_2 _10060_ (.A1(_01682_),
    .A2(_01684_),
    .B1(_02363_),
    .C1(_02364_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21oi_4 _10061_ (.A1(_02302_),
    .A2(_02366_),
    .B1(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__xnor2_4 _10062_ (.A(_03037_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__xnor2_4 _10063_ (.A(_02947_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__a21boi_4 _10064_ (.A1(_02264_),
    .A2(_02370_),
    .B1_N(_02369_),
    .Y(_03043_));
 sky130_fd_sc_hd__xor2_4 _10065_ (.A(_03041_),
    .B(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__xnor2_4 _10066_ (.A(_02890_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__a21bo_1 _10067_ (.A1(_02197_),
    .A2(_02375_),
    .B1_N(_02374_),
    .X(_03046_));
 sky130_fd_sc_hd__xnor2_4 _10068_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__xnor2_4 _10069_ (.A(_02793_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21boi_4 _10070_ (.A1(_02109_),
    .A2(_02379_),
    .B1_N(_02378_),
    .Y(_03049_));
 sky130_fd_sc_hd__xor2_4 _10071_ (.A(_03048_),
    .B(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__xnor2_4 _10072_ (.A(_02666_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__a21boi_2 _10073_ (.A1(_01973_),
    .A2(_02384_),
    .B1_N(_02382_),
    .Y(_03052_));
 sky130_fd_sc_hd__xor2_2 _10074_ (.A(_03051_),
    .B(_03052_),
    .X(_03054_));
 sky130_fd_sc_hd__xnor2_1 _10075_ (.A(_02451_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__a21boi_1 _10076_ (.A1(_01764_),
    .A2(_02388_),
    .B1_N(_02387_),
    .Y(_03056_));
 sky130_fd_sc_hd__xnor2_1 _10077_ (.A(_03055_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__xor2_1 _10078_ (.A(_02409_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__a21oi_1 _10079_ (.A1(_02391_),
    .A2(_02393_),
    .B1(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__and3_1 _10080_ (.A(_02391_),
    .B(_02393_),
    .C(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__nor2_1 _10081_ (.A(_03059_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__nand3b_1 _10082_ (.A_N(net286),
    .B(_01715_),
    .C(_01717_),
    .Y(_03062_));
 sky130_fd_sc_hd__o211ai_1 _10083_ (.A1(_01712_),
    .A2(net286),
    .B1(_02393_),
    .C1(_02395_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21oi_1 _10084_ (.A1(_03062_),
    .A2(_03063_),
    .B1(_02397_),
    .Y(_03064_));
 sky130_fd_sc_hd__a41o_4 _10085_ (.A1(_01132_),
    .A2(_01133_),
    .A3(_01718_),
    .A4(_02398_),
    .B1(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__xor2_1 _10086_ (.A(_03061_),
    .B(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__and2_1 _10087_ (.A(net284),
    .B(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__or2_1 _10088_ (.A(net284),
    .B(_03066_),
    .X(_03068_));
 sky130_fd_sc_hd__or2b_1 _10089_ (.A(_03067_),
    .B_N(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__inv_2 _10090_ (.A(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__a21o_1 _10091_ (.A1(_02403_),
    .A2(_02406_),
    .B1(_02402_),
    .X(_03071_));
 sky130_fd_sc_hd__a21oi_1 _10092_ (.A1(_03070_),
    .A2(_03071_),
    .B1(_00166_),
    .Y(_03072_));
 sky130_fd_sc_hd__o21a_1 _10093_ (.A1(_03070_),
    .A2(_03071_),
    .B1(_03072_),
    .X(_00008_));
 sky130_fd_sc_hd__a21o_1 _10094_ (.A1(_02391_),
    .A2(_02393_),
    .B1(_03058_),
    .X(_03074_));
 sky130_fd_sc_hd__a21bo_1 _10095_ (.A1(_03061_),
    .A2(_03065_),
    .B1_N(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__or2_1 _10096_ (.A(_03055_),
    .B(_03056_),
    .X(_03076_));
 sky130_fd_sc_hd__or2b_1 _10097_ (.A(_03057_),
    .B_N(_02409_),
    .X(_03077_));
 sky130_fd_sc_hd__or2b_1 _10098_ (.A(_02450_),
    .B_N(_02411_),
    .X(_03078_));
 sky130_fd_sc_hd__o21ai_2 _10099_ (.A1(_02412_),
    .A2(_02449_),
    .B1(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__and2b_1 _10100_ (.A_N(_02446_),
    .B(_02416_),
    .X(_03080_));
 sky130_fd_sc_hd__a21o_1 _10101_ (.A1(_02414_),
    .A2(_02447_),
    .B1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__a21o_2 _10102_ (.A1(_02453_),
    .A2(_02664_),
    .B1(_02663_),
    .X(_03082_));
 sky130_fd_sc_hd__or2b_1 _10103_ (.A(_02444_),
    .B_N(_02418_),
    .X(_03083_));
 sky130_fd_sc_hd__or2b_1 _10104_ (.A(_02445_),
    .B_N(_02417_),
    .X(_03085_));
 sky130_fd_sc_hd__nand2_2 _10105_ (.A(_03083_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__inv_2 _10106_ (.A(_02484_),
    .Y(_03087_));
 sky130_fd_sc_hd__or2b_1 _10107_ (.A(_02575_),
    .B_N(_02576_),
    .X(_03088_));
 sky130_fd_sc_hd__o21a_2 _10108_ (.A1(_03087_),
    .A2(_02577_),
    .B1(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__o21ba_2 _10109_ (.A1(_02438_),
    .A2(_02439_),
    .B1_N(_02443_),
    .X(_03090_));
 sky130_fd_sc_hd__or2b_1 _10110_ (.A(_02482_),
    .B_N(_02455_),
    .X(_03091_));
 sky130_fd_sc_hd__or2b_1 _10111_ (.A(_02454_),
    .B_N(_02483_),
    .X(_03092_));
 sky130_fd_sc_hd__or2b_1 _10112_ (.A(_02424_),
    .B_N(_02419_),
    .X(_03093_));
 sky130_fd_sc_hd__or2b_1 _10113_ (.A(_02427_),
    .B_N(_02425_),
    .X(_03094_));
 sky130_fd_sc_hd__a22o_1 _10114_ (.A1(net170),
    .A2(net162),
    .B1(_01188_),
    .B2(net169),
    .X(_03096_));
 sky130_fd_sc_hd__nand4_1 _10115_ (.A(net169),
    .B(_00171_),
    .C(_01777_),
    .D(_01188_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_03096_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__nand2_1 _10117_ (.A(_00270_),
    .B(net171),
    .Y(_03099_));
 sky130_fd_sc_hd__xor2_1 _10118_ (.A(_03098_),
    .B(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__xnor2_1 _10119_ (.A(_02466_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__o21ai_1 _10120_ (.A1(_02422_),
    .A2(_02423_),
    .B1(_02421_),
    .Y(_03102_));
 sky130_fd_sc_hd__xor2_1 _10121_ (.A(_03101_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__a21oi_1 _10122_ (.A1(_03093_),
    .A2(_03094_),
    .B1(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__and3_1 _10123_ (.A(_03093_),
    .B(_03094_),
    .C(_03103_),
    .X(_03105_));
 sky130_fd_sc_hd__nor2_1 _10124_ (.A(_03104_),
    .B(_03105_),
    .Y(_03107_));
 sky130_fd_sc_hd__and2_1 _10125_ (.A(_06243_),
    .B(net172),
    .X(_03108_));
 sky130_fd_sc_hd__nor2_1 _10126_ (.A(_03107_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__and2_1 _10127_ (.A(_03107_),
    .B(_03108_),
    .X(_03110_));
 sky130_fd_sc_hd__or2_1 _10128_ (.A(_03109_),
    .B(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__a21oi_1 _10129_ (.A1(_02431_),
    .A2(_02436_),
    .B1(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__and3_1 _10130_ (.A(_02431_),
    .B(_02436_),
    .C(_03111_),
    .X(_03113_));
 sky130_fd_sc_hd__nor2_1 _10131_ (.A(_03112_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__nand2_1 _10132_ (.A(_06127_),
    .B(net173),
    .Y(_03115_));
 sky130_fd_sc_hd__xor2_1 _10133_ (.A(_03114_),
    .B(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__a21oi_1 _10134_ (.A1(_03091_),
    .A2(_03092_),
    .B1(_03116_),
    .Y(_03118_));
 sky130_fd_sc_hd__and3_1 _10135_ (.A(_03091_),
    .B(_03092_),
    .C(_03116_),
    .X(_03119_));
 sky130_fd_sc_hd__nor2_2 _10136_ (.A(_03118_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__xnor2_4 _10137_ (.A(_03090_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_4 _10138_ (.A(_03089_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__xnor2_4 _10139_ (.A(_03086_),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__xor2_2 _10140_ (.A(_03082_),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__xnor2_2 _10141_ (.A(_03081_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__nand2_2 _10142_ (.A(_02659_),
    .B(_02661_),
    .Y(_03126_));
 sky130_fd_sc_hd__and2b_1 _10143_ (.A_N(_02791_),
    .B(_02669_),
    .X(_03127_));
 sky130_fd_sc_hd__a21o_2 _10144_ (.A1(_02667_),
    .A2(_02792_),
    .B1(_03127_),
    .X(_03129_));
 sky130_fd_sc_hd__or2b_1 _10145_ (.A(_02479_),
    .B_N(_02458_),
    .X(_03130_));
 sky130_fd_sc_hd__a21bo_2 _10146_ (.A1(_02457_),
    .A2(_02480_),
    .B1_N(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__nor2_2 _10147_ (.A(_02538_),
    .B(_02540_),
    .Y(_03132_));
 sky130_fd_sc_hd__or2b_1 _10148_ (.A(_02477_),
    .B_N(_02463_),
    .X(_03133_));
 sky130_fd_sc_hd__or2b_1 _10149_ (.A(_02478_),
    .B_N(_02461_),
    .X(_03134_));
 sky130_fd_sc_hd__nand2_4 _10150_ (.A(_03133_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_2 _10151_ (.A(_02511_),
    .B(_02513_),
    .Y(_03136_));
 sky130_fd_sc_hd__or2_1 _10152_ (.A(_02474_),
    .B(_02475_),
    .X(_03137_));
 sky130_fd_sc_hd__o21ai_2 _10153_ (.A1(_02467_),
    .A2(_02476_),
    .B1(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__and2b_1 _10154_ (.A_N(_02485_),
    .B(_02494_),
    .X(_03140_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_06130_),
    .B(_02464_),
    .Y(_03141_));
 sky130_fd_sc_hd__a22o_1 _10156_ (.A1(net19),
    .A2(net29),
    .B1(net30),
    .B2(net18),
    .X(_03142_));
 sky130_fd_sc_hd__nand4_1 _10157_ (.A(net18),
    .B(net19),
    .C(_00647_),
    .D(_01181_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_03142_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_1 _10159_ (.A(_06138_),
    .B(net31),
    .Y(_03145_));
 sky130_fd_sc_hd__xnor2_2 _10160_ (.A(_03144_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__or2_1 _10161_ (.A(_02471_),
    .B(_02473_),
    .X(_03147_));
 sky130_fd_sc_hd__xnor2_2 _10162_ (.A(_03146_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__xnor2_1 _10163_ (.A(_03141_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__o21a_1 _10164_ (.A1(_02491_),
    .A2(_03140_),
    .B1(_03149_),
    .X(_03151_));
 sky130_fd_sc_hd__nor3_1 _10165_ (.A(_02491_),
    .B(_03140_),
    .C(_03149_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor2_1 _10166_ (.A(_03151_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__xnor2_2 _10167_ (.A(_03138_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__xnor2_4 _10168_ (.A(_03136_),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__xor2_4 _10169_ (.A(_03135_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__xor2_4 _10170_ (.A(_03132_),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__xor2_4 _10171_ (.A(_03131_),
    .B(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__o21ai_1 _10172_ (.A1(_01886_),
    .A2(_01888_),
    .B1(_02572_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_02542_),
    .B(_02574_),
    .Y(_03160_));
 sky130_fd_sc_hd__a22o_1 _10174_ (.A1(net27),
    .A2(net21),
    .B1(net22),
    .B2(net26),
    .X(_03162_));
 sky130_fd_sc_hd__nand4_1 _10175_ (.A(net26),
    .B(net27),
    .C(net21),
    .D(net22),
    .Y(_03163_));
 sky130_fd_sc_hd__and2_1 _10176_ (.A(_03162_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(_00250_),
    .B(_00706_),
    .Y(_03165_));
 sky130_fd_sc_hd__xnor2_1 _10178_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__xnor2_1 _10179_ (.A(_02500_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21oi_1 _10180_ (.A1(_02488_),
    .A2(_02490_),
    .B1(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__and3_1 _10181_ (.A(_02488_),
    .B(_02490_),
    .C(_03167_),
    .X(_03169_));
 sky130_fd_sc_hd__nor2_1 _10182_ (.A(_03168_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__nor3_1 _10183_ (.A(_02499_),
    .B(_02500_),
    .C(_02509_),
    .Y(_03171_));
 sky130_fd_sc_hd__a22oi_1 _10184_ (.A1(_00238_),
    .A2(net91),
    .B1(net99),
    .B2(net90),
    .Y(_03173_));
 sky130_fd_sc_hd__and4_1 _10185_ (.A(net90),
    .B(net98),
    .C(net91),
    .D(net99),
    .X(_03174_));
 sky130_fd_sc_hd__o2bb2a_1 _10186_ (.A1_N(_06284_),
    .A2_N(net101),
    .B1(_03173_),
    .B2(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__and4bb_1 _10187_ (.A_N(_03173_),
    .B_N(_03174_),
    .C(net88),
    .D(net101),
    .X(_03176_));
 sky130_fd_sc_hd__or2_1 _10188_ (.A(_03175_),
    .B(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__nand2_1 _10189_ (.A(_02504_),
    .B(_02506_),
    .Y(_03178_));
 sky130_fd_sc_hd__xnor2_1 _10190_ (.A(_03177_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__clkbuf_4 _10191_ (.A(net102),
    .X(_03180_));
 sky130_fd_sc_hd__nand2_1 _10192_ (.A(_06159_),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__xnor2_1 _10193_ (.A(_03179_),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__o21a_1 _10194_ (.A1(_02507_),
    .A2(_03171_),
    .B1(_03182_),
    .X(_03184_));
 sky130_fd_sc_hd__nor3_1 _10195_ (.A(_02507_),
    .B(_03171_),
    .C(_03182_),
    .Y(_03185_));
 sky130_fd_sc_hd__nor2_1 _10196_ (.A(_03184_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__xnor2_1 _10197_ (.A(_03170_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__a21bo_1 _10198_ (.A1(_02522_),
    .A2(_02530_),
    .B1_N(_02529_),
    .X(_03188_));
 sky130_fd_sc_hd__and3b_1 _10199_ (.A_N(_02555_),
    .B(_02556_),
    .C(_02548_),
    .X(_03189_));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_02526_),
    .B(_02528_),
    .Y(_03190_));
 sky130_fd_sc_hd__nand2_1 _10201_ (.A(_06254_),
    .B(net93),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _10202_ (.A(net97),
    .B(net92),
    .Y(_03192_));
 sky130_fd_sc_hd__xor2_1 _10203_ (.A(_03191_),
    .B(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__xor2_1 _10204_ (.A(_02546_),
    .B(_03193_),
    .X(_03195_));
 sky130_fd_sc_hd__xor2_1 _10205_ (.A(_03190_),
    .B(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__o21a_1 _10206_ (.A1(_02555_),
    .A2(_03189_),
    .B1(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__or3_1 _10207_ (.A(_02555_),
    .B(_03189_),
    .C(_03196_),
    .X(_03198_));
 sky130_fd_sc_hd__and2b_1 _10208_ (.A_N(_03197_),
    .B(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__xnor2_1 _10209_ (.A(_03188_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o21ba_1 _10210_ (.A1(_02520_),
    .A2(_02534_),
    .B1_N(_02533_),
    .X(_03201_));
 sky130_fd_sc_hd__xor2_1 _10211_ (.A(_03200_),
    .B(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__xnor2_1 _10212_ (.A(_03187_),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__and2b_1 _10213_ (.A_N(_02566_),
    .B(_02567_),
    .X(_03204_));
 sky130_fd_sc_hd__or2b_1 _10214_ (.A(_02567_),
    .B_N(_02566_),
    .X(_03206_));
 sky130_fd_sc_hd__o21ai_2 _10215_ (.A1(_02559_),
    .A2(_03204_),
    .B1(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _10216_ (.A(_01947_),
    .B(_01949_),
    .Y(_03208_));
 sky130_fd_sc_hd__a21oi_2 _10217_ (.A1(_03208_),
    .A2(_02607_),
    .B1(_02606_),
    .Y(_03209_));
 sky130_fd_sc_hd__clkbuf_4 _10218_ (.A(net138),
    .X(_03210_));
 sky130_fd_sc_hd__a22oi_1 _10219_ (.A1(_06274_),
    .A2(_01250_),
    .B1(_03210_),
    .B2(_06152_),
    .Y(_03211_));
 sky130_fd_sc_hd__and4_2 _10220_ (.A(_06152_),
    .B(_06274_),
    .C(_01250_),
    .D(_03210_),
    .X(_03212_));
 sky130_fd_sc_hd__nor2_2 _10221_ (.A(_03211_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__and4_1 _10222_ (.A(_06283_),
    .B(_00210_),
    .C(_00201_),
    .D(_00677_),
    .X(_03214_));
 sky130_fd_sc_hd__and4_1 _10223_ (.A(_06274_),
    .B(_00665_),
    .C(_02551_),
    .D(_02552_),
    .X(_03215_));
 sky130_fd_sc_hd__a22o_1 _10224_ (.A1(net135),
    .A2(net127),
    .B1(net128),
    .B2(net133),
    .X(_03217_));
 sky130_fd_sc_hd__nand4_1 _10225_ (.A(_06283_),
    .B(_00201_),
    .C(_00677_),
    .D(net128),
    .Y(_03218_));
 sky130_fd_sc_hd__and2_1 _10226_ (.A(net126),
    .B(net136),
    .X(_03219_));
 sky130_fd_sc_hd__a21o_1 _10227_ (.A1(_03217_),
    .A2(_03218_),
    .B1(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__nand3_1 _10228_ (.A(_03217_),
    .B(_03218_),
    .C(_03219_),
    .Y(_03221_));
 sky130_fd_sc_hd__o211ai_1 _10229_ (.A1(_03214_),
    .A2(_03215_),
    .B1(_03220_),
    .C1(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__a211o_1 _10230_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03214_),
    .C1(_03215_),
    .X(_03223_));
 sky130_fd_sc_hd__nand2_1 _10231_ (.A(_03222_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__xor2_2 _10232_ (.A(_03213_),
    .B(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__and2_1 _10233_ (.A(_02561_),
    .B(_02564_),
    .X(_03226_));
 sky130_fd_sc_hd__a21o_1 _10234_ (.A1(_02560_),
    .A2(_02565_),
    .B1(_03226_),
    .X(_03228_));
 sky130_fd_sc_hd__and4_1 _10235_ (.A(_06177_),
    .B(net142),
    .C(net153),
    .D(net154),
    .X(_03229_));
 sky130_fd_sc_hd__a31o_1 _10236_ (.A1(_04128_),
    .A2(net155),
    .A3(_02589_),
    .B1(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__nand2_1 _10237_ (.A(_04314_),
    .B(_01264_),
    .Y(_03231_));
 sky130_fd_sc_hd__and3_1 _10238_ (.A(_06151_),
    .B(_01872_),
    .C(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__xor2_2 _10239_ (.A(_03230_),
    .B(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__xor2_1 _10240_ (.A(_03228_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__xnor2_2 _10241_ (.A(_03225_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__xnor2_2 _10242_ (.A(_03209_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__xnor2_2 _10243_ (.A(_03207_),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__and2_1 _10244_ (.A(_02544_),
    .B(_02570_),
    .X(_03239_));
 sky130_fd_sc_hd__a21oi_2 _10245_ (.A1(_02543_),
    .A2(_02571_),
    .B1(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__xor2_1 _10246_ (.A(_03237_),
    .B(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__and2_1 _10247_ (.A(_03203_),
    .B(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__nor2_1 _10248_ (.A(_03203_),
    .B(_03241_),
    .Y(_03243_));
 sky130_fd_sc_hd__or2_1 _10249_ (.A(_03242_),
    .B(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__a21oi_1 _10250_ (.A1(_03159_),
    .A2(_03160_),
    .B1(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__and3_1 _10251_ (.A(_03159_),
    .B(_03160_),
    .C(_03244_),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_2 _10252_ (.A(_03245_),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__xnor2_4 _10253_ (.A(_03158_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__or2_1 _10254_ (.A(_02650_),
    .B(_02652_),
    .X(_03250_));
 sky130_fd_sc_hd__or2_1 _10255_ (.A(_02744_),
    .B(_02747_),
    .X(_03251_));
 sky130_fd_sc_hd__o21a_1 _10256_ (.A1(_02687_),
    .A2(_02748_),
    .B1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__nand2_1 _10257_ (.A(_02645_),
    .B(_02648_),
    .Y(_03253_));
 sky130_fd_sc_hd__a21o_1 _10258_ (.A1(_02670_),
    .A2(_02685_),
    .B1(_02684_),
    .X(_03254_));
 sky130_fd_sc_hd__nand2_2 _10259_ (.A(_02601_),
    .B(_02604_),
    .Y(_03255_));
 sky130_fd_sc_hd__a21o_1 _10260_ (.A1(_02612_),
    .A2(_02619_),
    .B1(_02618_),
    .X(_03256_));
 sky130_fd_sc_hd__and3_1 _10261_ (.A(net142),
    .B(net143),
    .C(net154),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _10262_ (.A1(_00291_),
    .A2(net153),
    .B1(_01288_),
    .B2(net142),
    .X(_03258_));
 sky130_fd_sc_hd__a21bo_1 _10263_ (.A1(_00749_),
    .A2(_03257_),
    .B1_N(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(_06178_),
    .B(net155),
    .Y(_03261_));
 sky130_fd_sc_hd__xor2_1 _10265_ (.A(_03259_),
    .B(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__a22o_1 _10266_ (.A1(net151),
    .A2(net146),
    .B1(net147),
    .B2(net150),
    .X(_03263_));
 sky130_fd_sc_hd__nand4_1 _10267_ (.A(_06171_),
    .B(_06319_),
    .C(net146),
    .D(net147),
    .Y(_03264_));
 sky130_fd_sc_hd__and2_1 _10268_ (.A(_01293_),
    .B(net144),
    .X(_03265_));
 sky130_fd_sc_hd__a21o_1 _10269_ (.A1(_03263_),
    .A2(_03264_),
    .B1(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__nand3_1 _10270_ (.A(_03263_),
    .B(_03264_),
    .C(_03265_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21bo_1 _10271_ (.A1(_02596_),
    .A2(_02598_),
    .B1_N(_02597_),
    .X(_03268_));
 sky130_fd_sc_hd__nand3_1 _10272_ (.A(_03266_),
    .B(_03267_),
    .C(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__a21o_1 _10273_ (.A1(_03266_),
    .A2(_03267_),
    .B1(_03268_),
    .X(_03270_));
 sky130_fd_sc_hd__nand3_1 _10274_ (.A(_03262_),
    .B(_03269_),
    .C(_03270_),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_1 _10275_ (.A1(_03269_),
    .A2(_03270_),
    .B1(_03262_),
    .X(_03273_));
 sky130_fd_sc_hd__and3_1 _10276_ (.A(_03256_),
    .B(_03272_),
    .C(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__a21o_1 _10277_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03256_),
    .X(_03275_));
 sky130_fd_sc_hd__or2b_1 _10278_ (.A(_03274_),
    .B_N(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__xnor2_2 _10279_ (.A(_03255_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__and4_1 _10280_ (.A(_06361_),
    .B(net204),
    .C(net213),
    .D(net214),
    .X(_03278_));
 sky130_fd_sc_hd__a31o_1 _10281_ (.A1(_06086_),
    .A2(net215),
    .A3(_02623_),
    .B1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_06086_),
    .B(net216),
    .Y(_03280_));
 sky130_fd_sc_hd__xor2_1 _10283_ (.A(_03279_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__and2_1 _10284_ (.A(_02616_),
    .B(_03281_),
    .X(_03283_));
 sky130_fd_sc_hd__nor2_1 _10285_ (.A(_02616_),
    .B(_03281_),
    .Y(_03284_));
 sky130_fd_sc_hd__or2_1 _10286_ (.A(_03283_),
    .B(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__a22oi_1 _10287_ (.A1(_00297_),
    .A2(_00810_),
    .B1(_00757_),
    .B2(_00343_),
    .Y(_03286_));
 sky130_fd_sc_hd__and4_1 _10288_ (.A(_00343_),
    .B(net213),
    .C(net205),
    .D(net214),
    .X(_03287_));
 sky130_fd_sc_hd__nor2_1 _10289_ (.A(_03286_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__nand2_1 _10290_ (.A(_06362_),
    .B(_02626_),
    .Y(_03289_));
 sky130_fd_sc_hd__xnor2_2 _10291_ (.A(_03288_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__a22oi_1 _10292_ (.A1(_06304_),
    .A2(_01365_),
    .B1(_01986_),
    .B2(_06173_),
    .Y(_03291_));
 sky130_fd_sc_hd__and4_1 _10293_ (.A(_06173_),
    .B(_06304_),
    .C(net206),
    .D(net207),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_1 _10294_ (.A(_03291_),
    .B(_03292_),
    .Y(_03294_));
 sky130_fd_sc_hd__a21bo_1 _10295_ (.A1(_02629_),
    .A2(_02631_),
    .B1_N(_02630_),
    .X(_03295_));
 sky130_fd_sc_hd__xor2_2 _10296_ (.A(_03294_),
    .B(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__xor2_2 _10297_ (.A(_03290_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__a21bo_1 _10298_ (.A1(_02628_),
    .A2(_02637_),
    .B1_N(_02636_),
    .X(_03298_));
 sky130_fd_sc_hd__xor2_1 _10299_ (.A(_03297_),
    .B(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__xnor2_2 _10300_ (.A(_03285_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__o21ba_1 _10301_ (.A1(_02621_),
    .A2(_02642_),
    .B1_N(_02641_),
    .X(_03301_));
 sky130_fd_sc_hd__xnor2_2 _10302_ (.A(_03300_),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__xor2_2 _10303_ (.A(_03277_),
    .B(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_2 _10304_ (.A(_03254_),
    .B(_03303_),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_2 _10305_ (.A(_03253_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_2 _10306_ (.A(_03252_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__xnor2_1 _10307_ (.A(_03250_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__a21boi_1 _10308_ (.A1(_02581_),
    .A2(_02655_),
    .B1_N(_02654_),
    .Y(_03309_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__and2_1 _10310_ (.A(_03308_),
    .B(_03309_),
    .X(_03311_));
 sky130_fd_sc_hd__nor2_2 _10311_ (.A(_03310_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__xnor2_4 _10312_ (.A(_03248_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__xnor2_4 _10313_ (.A(_03129_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__xor2_4 _10314_ (.A(_03126_),
    .B(_03314_),
    .X(_03316_));
 sky130_fd_sc_hd__a21o_2 _10315_ (.A1(_02749_),
    .A2(_02788_),
    .B1(_02787_),
    .X(_03317_));
 sky130_fd_sc_hd__a21o_1 _10316_ (.A1(_02795_),
    .A2(_02887_),
    .B1(_02886_),
    .X(_03318_));
 sky130_fd_sc_hd__or2b_1 _10317_ (.A(_02680_),
    .B_N(_02672_),
    .X(_03319_));
 sky130_fd_sc_hd__a21bo_2 _10318_ (.A1(_02671_),
    .A2(_02681_),
    .B1_N(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__a21bo_2 _10319_ (.A1(_02704_),
    .A2(_02719_),
    .B1_N(_02718_),
    .X(_03321_));
 sky130_fd_sc_hd__nor2_1 _10320_ (.A(_02674_),
    .B(_02677_),
    .Y(_03322_));
 sky130_fd_sc_hd__a21o_2 _10321_ (.A1(_02673_),
    .A2(_02678_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__a21oi_4 _10322_ (.A1(_02693_),
    .A2(_02702_),
    .B1(_02700_),
    .Y(_03324_));
 sky130_fd_sc_hd__a32oi_4 _10323_ (.A1(_06384_),
    .A2(net249),
    .A3(_02689_),
    .B1(_02688_),
    .B2(_01385_),
    .Y(_03325_));
 sky130_fd_sc_hd__a22o_1 _10324_ (.A1(_06384_),
    .A2(net250),
    .B1(_01987_),
    .B2(net237),
    .X(_03327_));
 sky130_fd_sc_hd__nand4_4 _10325_ (.A(net237),
    .B(net238),
    .C(net250),
    .D(net251),
    .Y(_03328_));
 sky130_fd_sc_hd__nand2_2 _10326_ (.A(_03327_),
    .B(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__xor2_4 _10327_ (.A(_03325_),
    .B(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__xnor2_4 _10328_ (.A(_02676_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__xor2_4 _10329_ (.A(_03324_),
    .B(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__xnor2_4 _10330_ (.A(_03323_),
    .B(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__xnor2_4 _10331_ (.A(_03321_),
    .B(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__xnor2_4 _10332_ (.A(_03320_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__a22o_1 _10333_ (.A1(net248),
    .A2(net240),
    .B1(net241),
    .B2(net247),
    .X(_03336_));
 sky130_fd_sc_hd__nand4_1 _10334_ (.A(net247),
    .B(net248),
    .C(net240),
    .D(net241),
    .Y(_03338_));
 sky130_fd_sc_hd__and2_1 _10335_ (.A(net239),
    .B(net249),
    .X(_03339_));
 sky130_fd_sc_hd__a21o_1 _10336_ (.A1(_03336_),
    .A2(_03338_),
    .B1(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__nand3_1 _10337_ (.A(_03336_),
    .B(_03338_),
    .C(_03339_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_2 _10338_ (.A(_03340_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand2_1 _10339_ (.A(_03864_),
    .B(_02694_),
    .Y(_03343_));
 sky130_fd_sc_hd__and3_2 _10340_ (.A(_05969_),
    .B(_02695_),
    .C(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__xnor2_4 _10341_ (.A(_03342_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__nand2_1 _10342_ (.A(_02708_),
    .B(_02710_),
    .Y(_03346_));
 sky130_fd_sc_hd__a22o_1 _10343_ (.A1(net2),
    .A2(net11),
    .B1(net13),
    .B2(net255),
    .X(_03347_));
 sky130_fd_sc_hd__nand4_1 _10344_ (.A(_06375_),
    .B(_00357_),
    .C(net11),
    .D(net13),
    .Y(_03349_));
 sky130_fd_sc_hd__and2_1 _10345_ (.A(net254),
    .B(net14),
    .X(_03350_));
 sky130_fd_sc_hd__a21oi_1 _10346_ (.A1(_03347_),
    .A2(_03349_),
    .B1(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__and3_1 _10347_ (.A(_03347_),
    .B(_03349_),
    .C(_03350_),
    .X(_03352_));
 sky130_fd_sc_hd__a211o_1 _10348_ (.A1(_02727_),
    .A2(_02729_),
    .B1(_03351_),
    .C1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__o211ai_2 _10349_ (.A1(_03351_),
    .A2(_03352_),
    .B1(_02727_),
    .C1(_02729_),
    .Y(_03354_));
 sky130_fd_sc_hd__nand3_1 _10350_ (.A(_03346_),
    .B(_03353_),
    .C(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21o_1 _10351_ (.A1(_03353_),
    .A2(_03354_),
    .B1(_03346_),
    .X(_03356_));
 sky130_fd_sc_hd__a21bo_1 _10352_ (.A1(_02705_),
    .A2(_02713_),
    .B1_N(_02711_),
    .X(_03357_));
 sky130_fd_sc_hd__and3_1 _10353_ (.A(_03355_),
    .B(_03356_),
    .C(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__a21o_1 _10354_ (.A1(_03355_),
    .A2(_03356_),
    .B1(_03357_),
    .X(_03360_));
 sky130_fd_sc_hd__or2b_2 _10355_ (.A(_03358_),
    .B_N(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__xnor2_4 _10356_ (.A(_03345_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__nor3_1 _10357_ (.A(_02732_),
    .B(_02733_),
    .C(_02736_),
    .Y(_03363_));
 sky130_fd_sc_hd__a31o_1 _10358_ (.A1(_02728_),
    .A2(_02729_),
    .A3(_02737_),
    .B1(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__a21o_1 _10359_ (.A1(_02754_),
    .A2(_02762_),
    .B1(_02761_),
    .X(_03365_));
 sky130_fd_sc_hd__a22oi_1 _10360_ (.A1(_06368_),
    .A2(net4),
    .B1(net5),
    .B2(_05882_),
    .Y(_03366_));
 sky130_fd_sc_hd__and4_1 _10361_ (.A(net8),
    .B(net9),
    .C(net4),
    .D(net5),
    .X(_03367_));
 sky130_fd_sc_hd__nor2_1 _10362_ (.A(_03366_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(net10),
    .B(_00850_),
    .Y(_03369_));
 sky130_fd_sc_hd__xnor2_2 _10364_ (.A(_03368_),
    .B(_03369_),
    .Y(_03371_));
 sky130_fd_sc_hd__a21o_1 _10365_ (.A1(_05750_),
    .A2(net66),
    .B1(_02733_),
    .X(_03372_));
 sky130_fd_sc_hd__a21bo_1 _10366_ (.A1(_05750_),
    .A2(_02733_),
    .B1_N(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__xnor2_2 _10367_ (.A(_03371_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__xor2_2 _10368_ (.A(_03365_),
    .B(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__xor2_2 _10369_ (.A(_03364_),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__and2b_1 _10370_ (.A_N(_02725_),
    .B(_02738_),
    .X(_03377_));
 sky130_fd_sc_hd__a21o_1 _10371_ (.A1(_02724_),
    .A2(_02739_),
    .B1(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__xor2_2 _10372_ (.A(_03376_),
    .B(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__xnor2_2 _10373_ (.A(_03362_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__and2b_1 _10374_ (.A_N(_02742_),
    .B(_02740_),
    .X(_03382_));
 sky130_fd_sc_hd__a21oi_2 _10375_ (.A1(_02722_),
    .A2(_02743_),
    .B1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__xnor2_2 _10376_ (.A(_03380_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_2 _10377_ (.A(_03335_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__or2b_1 _10378_ (.A(_02753_),
    .B_N(_02781_),
    .X(_03386_));
 sky130_fd_sc_hd__a21bo_1 _10379_ (.A1(_02752_),
    .A2(_02782_),
    .B1_N(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__a21oi_2 _10380_ (.A1(_02814_),
    .A2(_02850_),
    .B1(_02848_),
    .Y(_03388_));
 sky130_fd_sc_hd__or2b_1 _10381_ (.A(_02779_),
    .B_N(_02777_),
    .X(_03389_));
 sky130_fd_sc_hd__or2b_1 _10382_ (.A(_02764_),
    .B_N(_02780_),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_03389_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__a21o_1 _10384_ (.A1(_02796_),
    .A2(_02812_),
    .B1(_02810_),
    .X(_03393_));
 sky130_fd_sc_hd__nand2_2 _10385_ (.A(_02758_),
    .B(_02760_),
    .Y(_03394_));
 sky130_fd_sc_hd__a32o_1 _10386_ (.A1(_06347_),
    .A2(_00879_),
    .A3(_02768_),
    .B1(_02766_),
    .B2(_02765_),
    .X(_03395_));
 sky130_fd_sc_hd__a22o_1 _10387_ (.A1(net63),
    .A2(net55),
    .B1(net64),
    .B2(net54),
    .X(_03396_));
 sky130_fd_sc_hd__nand4_2 _10388_ (.A(net54),
    .B(net63),
    .C(net55),
    .D(net64),
    .Y(_03397_));
 sky130_fd_sc_hd__a22o_1 _10389_ (.A1(_06343_),
    .A2(net65),
    .B1(_03396_),
    .B2(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__nand4_2 _10390_ (.A(_06343_),
    .B(net65),
    .C(_03396_),
    .D(_03397_),
    .Y(_03399_));
 sky130_fd_sc_hd__and3_1 _10391_ (.A(_03395_),
    .B(_03398_),
    .C(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__a21o_1 _10392_ (.A1(_03398_),
    .A2(_03399_),
    .B1(_03395_),
    .X(_03401_));
 sky130_fd_sc_hd__and2b_1 _10393_ (.A_N(_03400_),
    .B(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__xnor2_2 _10394_ (.A(_03394_),
    .B(_03402_),
    .Y(_03404_));
 sky130_fd_sc_hd__a22oi_1 _10395_ (.A1(_06347_),
    .A2(_01444_),
    .B1(_02765_),
    .B2(_05761_),
    .Y(_03405_));
 sky130_fd_sc_hd__and4_1 _10396_ (.A(_05761_),
    .B(net62),
    .C(net57),
    .D(net58),
    .X(_03406_));
 sky130_fd_sc_hd__nor2_1 _10397_ (.A(_03405_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__a22o_1 _10398_ (.A1(_06424_),
    .A2(_01443_),
    .B1(_02064_),
    .B2(_05498_),
    .X(_03408_));
 sky130_fd_sc_hd__nand4_2 _10399_ (.A(net70),
    .B(net71),
    .C(net83),
    .D(net84),
    .Y(_03409_));
 sky130_fd_sc_hd__xor2_1 _10400_ (.A(_02773_),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__nand2_1 _10401_ (.A(_03408_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__xor2_2 _10402_ (.A(_03407_),
    .B(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__nor2_1 _10403_ (.A(_02774_),
    .B(_02775_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _10404_ (.A(_02774_),
    .B(_02775_),
    .Y(_03415_));
 sky130_fd_sc_hd__o21a_1 _10405_ (.A1(_02771_),
    .A2(_03413_),
    .B1(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__xnor2_2 _10406_ (.A(_03412_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__xor2_2 _10407_ (.A(_03404_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__xnor2_2 _10408_ (.A(_03393_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_2 _10409_ (.A(_03391_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__xnor2_2 _10410_ (.A(_03388_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__xnor2_2 _10411_ (.A(_03387_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__nor2_1 _10412_ (.A(_02751_),
    .B(_02783_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_2 _10413_ (.A1(_02750_),
    .A2(_02784_),
    .B1(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__xor2_1 _10414_ (.A(_03422_),
    .B(_03424_),
    .X(_03426_));
 sky130_fd_sc_hd__xnor2_1 _10415_ (.A(_03385_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__and2_1 _10416_ (.A(_03318_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__nor2_1 _10417_ (.A(_03318_),
    .B(_03427_),
    .Y(_03429_));
 sky130_fd_sc_hd__nor2_2 _10418_ (.A(_03428_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__xor2_4 _10419_ (.A(_03317_),
    .B(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_1 _10420_ (.A(_02882_),
    .B(_02884_),
    .Y(_03432_));
 sky130_fd_sc_hd__and2_1 _10421_ (.A(_02891_),
    .B(_02942_),
    .X(_03433_));
 sky130_fd_sc_hd__nand2_1 _10422_ (.A(_02806_),
    .B(_02808_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21o_1 _10423_ (.A1(_02818_),
    .A2(_02827_),
    .B1(_02826_),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_1 _10424_ (.A(_02803_),
    .B(_02805_),
    .Y(_03437_));
 sky130_fd_sc_hd__a22o_1 _10425_ (.A1(net81),
    .A2(net73),
    .B1(net74),
    .B2(net80),
    .X(_03438_));
 sky130_fd_sc_hd__nand4_1 _10426_ (.A(_06410_),
    .B(net81),
    .C(net73),
    .D(net74),
    .Y(_03439_));
 sky130_fd_sc_hd__a22o_1 _10427_ (.A1(_00431_),
    .A2(net82),
    .B1(_03438_),
    .B2(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__nand4_1 _10428_ (.A(_00431_),
    .B(net82),
    .C(_03438_),
    .D(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand3_1 _10429_ (.A(_02817_),
    .B(_03440_),
    .C(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__a21o_1 _10430_ (.A1(_03440_),
    .A2(_03441_),
    .B1(_02817_),
    .X(_03443_));
 sky130_fd_sc_hd__nand3_1 _10431_ (.A(_03437_),
    .B(_03442_),
    .C(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__a21o_1 _10432_ (.A1(_03442_),
    .A2(_03443_),
    .B1(_03437_),
    .X(_03445_));
 sky130_fd_sc_hd__and3_1 _10433_ (.A(_03435_),
    .B(_03444_),
    .C(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__a21o_1 _10434_ (.A1(_03444_),
    .A2(_03445_),
    .B1(_03435_),
    .X(_03448_));
 sky130_fd_sc_hd__or2b_1 _10435_ (.A(_03446_),
    .B_N(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__xnor2_1 _10436_ (.A(_03434_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__nand3_1 _10437_ (.A(_02840_),
    .B(_02841_),
    .C(_02842_),
    .Y(_03451_));
 sky130_fd_sc_hd__a21bo_1 _10438_ (.A1(_02832_),
    .A2(_02835_),
    .B1_N(_02834_),
    .X(_03452_));
 sky130_fd_sc_hd__inv_2 _10439_ (.A(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a22o_1 _10440_ (.A1(net116),
    .A2(net109),
    .B1(net110),
    .B2(net115),
    .X(_03454_));
 sky130_fd_sc_hd__nand4_1 _10441_ (.A(net115),
    .B(net116),
    .C(net109),
    .D(net110),
    .Y(_03455_));
 sky130_fd_sc_hd__a22o_1 _10442_ (.A1(net117),
    .A2(net108),
    .B1(_03454_),
    .B2(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nand4_1 _10443_ (.A(_00438_),
    .B(_00956_),
    .C(_03454_),
    .D(_03455_),
    .Y(_03457_));
 sky130_fd_sc_hd__and3_1 _10444_ (.A(_02859_),
    .B(_03456_),
    .C(_03457_),
    .X(_03459_));
 sky130_fd_sc_hd__a21oi_1 _10445_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_02859_),
    .Y(_03460_));
 sky130_fd_sc_hd__or3_1 _10446_ (.A(_03453_),
    .B(_03459_),
    .C(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__o21ai_1 _10447_ (.A1(_03459_),
    .A2(_03460_),
    .B1(_03453_),
    .Y(_03462_));
 sky130_fd_sc_hd__a21bo_1 _10448_ (.A1(_02830_),
    .A2(_02839_),
    .B1_N(_02838_),
    .X(_03463_));
 sky130_fd_sc_hd__and3_1 _10449_ (.A(_03461_),
    .B(_03462_),
    .C(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__a21o_1 _10450_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03463_),
    .X(_03465_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_05520_),
    .B(_02799_),
    .Y(_03466_));
 sky130_fd_sc_hd__a22o_1 _10452_ (.A1(net107),
    .A2(net118),
    .B1(net119),
    .B2(net106),
    .X(_03467_));
 sky130_fd_sc_hd__nand4_1 _10453_ (.A(_06437_),
    .B(_00454_),
    .C(net118),
    .D(net119),
    .Y(_03468_));
 sky130_fd_sc_hd__and2_1 _10454_ (.A(net105),
    .B(net120),
    .X(_03470_));
 sky130_fd_sc_hd__a21oi_1 _10455_ (.A1(_03467_),
    .A2(_03468_),
    .B1(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__and3_1 _10456_ (.A(_03467_),
    .B(_03468_),
    .C(_03470_),
    .X(_03472_));
 sky130_fd_sc_hd__a211oi_1 _10457_ (.A1(_02823_),
    .A2(_02825_),
    .B1(_03471_),
    .C1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__o211a_1 _10458_ (.A1(_03471_),
    .A2(_03472_),
    .B1(_02823_),
    .C1(_02825_),
    .X(_03474_));
 sky130_fd_sc_hd__nor2_1 _10459_ (.A(_03473_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__xnor2_1 _10460_ (.A(_03466_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__and3b_1 _10461_ (.A_N(_03464_),
    .B(_03465_),
    .C(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__a21oi_1 _10462_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03463_),
    .Y(_03478_));
 sky130_fd_sc_hd__o21ba_1 _10463_ (.A1(_03464_),
    .A2(_03478_),
    .B1_N(_03476_),
    .X(_03479_));
 sky130_fd_sc_hd__a211o_1 _10464_ (.A1(_03451_),
    .A2(_02846_),
    .B1(_03477_),
    .C1(_03479_),
    .X(_03481_));
 sky130_fd_sc_hd__o211ai_2 _10465_ (.A1(_03477_),
    .A2(_03479_),
    .B1(_03451_),
    .C1(_02846_),
    .Y(_03482_));
 sky130_fd_sc_hd__and3_1 _10466_ (.A(_03450_),
    .B(_03481_),
    .C(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__a21oi_1 _10467_ (.A1(_03481_),
    .A2(_03482_),
    .B1(_03450_),
    .Y(_03484_));
 sky130_fd_sc_hd__or2_2 _10468_ (.A(_03483_),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__nand3_1 _10469_ (.A(_02854_),
    .B(_02878_),
    .C(_02879_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(_02869_),
    .B(_02871_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21bo_1 _10471_ (.A1(_02892_),
    .A2(_02900_),
    .B1_N(_02898_),
    .X(_03488_));
 sky130_fd_sc_hd__a22o_1 _10472_ (.A1(net177),
    .A2(net134),
    .B1(net178),
    .B2(net123),
    .X(_03489_));
 sky130_fd_sc_hd__nand4_2 _10473_ (.A(_00479_),
    .B(net177),
    .C(net134),
    .D(net178),
    .Y(_03490_));
 sky130_fd_sc_hd__and2_1 _10474_ (.A(net111),
    .B(net180),
    .X(_03492_));
 sky130_fd_sc_hd__a21o_1 _10475_ (.A1(_03489_),
    .A2(_03490_),
    .B1(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__nand3_1 _10476_ (.A(_03489_),
    .B(_03490_),
    .C(_03492_),
    .Y(_03494_));
 sky130_fd_sc_hd__a21bo_1 _10477_ (.A1(_02863_),
    .A2(_02865_),
    .B1_N(_02864_),
    .X(_03495_));
 sky130_fd_sc_hd__nand3_1 _10478_ (.A(_03493_),
    .B(_03494_),
    .C(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__a21o_1 _10479_ (.A1(_03493_),
    .A2(_03494_),
    .B1(_03495_),
    .X(_03497_));
 sky130_fd_sc_hd__a22o_1 _10480_ (.A1(_05191_),
    .A2(net181),
    .B1(_03496_),
    .B2(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_4 _10481_ (.A(net181),
    .X(_03499_));
 sky130_fd_sc_hd__nand4_2 _10482_ (.A(_05191_),
    .B(_03499_),
    .C(_03496_),
    .D(_03497_),
    .Y(_03500_));
 sky130_fd_sc_hd__nand3_2 _10483_ (.A(_03488_),
    .B(_03498_),
    .C(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__a21o_1 _10484_ (.A1(_03498_),
    .A2(_03500_),
    .B1(_03488_),
    .X(_03503_));
 sky130_fd_sc_hd__and3_1 _10485_ (.A(_03487_),
    .B(_03501_),
    .C(_03503_),
    .X(_03504_));
 sky130_fd_sc_hd__a21oi_2 _10486_ (.A1(_03501_),
    .A2(_03503_),
    .B1(_03487_),
    .Y(_03505_));
 sky130_fd_sc_hd__a211oi_4 _10487_ (.A1(_02920_),
    .A2(_02923_),
    .B1(_03504_),
    .C1(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__o211a_1 _10488_ (.A1(_03504_),
    .A2(_03505_),
    .B1(_02920_),
    .C1(_02923_),
    .X(_03507_));
 sky130_fd_sc_hd__a211oi_4 _10489_ (.A1(_02873_),
    .A2(_02875_),
    .B1(_03506_),
    .C1(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__o211a_1 _10490_ (.A1(_03506_),
    .A2(_03507_),
    .B1(_02873_),
    .C1(_02875_),
    .X(_03509_));
 sky130_fd_sc_hd__a211oi_2 _10491_ (.A1(_02878_),
    .A2(_03486_),
    .B1(_03508_),
    .C1(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__o211a_1 _10492_ (.A1(_03508_),
    .A2(_03509_),
    .B1(_02878_),
    .C1(_03486_),
    .X(_03511_));
 sky130_fd_sc_hd__or3_1 _10493_ (.A(_03485_),
    .B(_03510_),
    .C(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__o21ai_1 _10494_ (.A1(_03510_),
    .A2(_03511_),
    .B1(_03485_),
    .Y(_03514_));
 sky130_fd_sc_hd__o211ai_2 _10495_ (.A1(_03433_),
    .A2(_02945_),
    .B1(_03512_),
    .C1(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a211o_1 _10496_ (.A1(_03512_),
    .A2(_03514_),
    .B1(_03433_),
    .C1(_02945_),
    .X(_03516_));
 sky130_fd_sc_hd__and3_1 _10497_ (.A(_03432_),
    .B(_03515_),
    .C(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__a21oi_1 _10498_ (.A1(_03515_),
    .A2(_03516_),
    .B1(_03432_),
    .Y(_03518_));
 sky130_fd_sc_hd__nor2_2 _10499_ (.A(_03517_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__or2b_1 _10500_ (.A(_02940_),
    .B_N(_02939_),
    .X(_03520_));
 sky130_fd_sc_hd__o21ai_4 _10501_ (.A1(_02925_),
    .A2(_02941_),
    .B1(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__and2b_1 _10502_ (.A_N(_02977_),
    .B(_02949_),
    .X(_03522_));
 sky130_fd_sc_hd__a21o_1 _10503_ (.A1(_02948_),
    .A2(_02978_),
    .B1(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__or2b_2 _10504_ (.A(_02895_),
    .B_N(_02897_),
    .X(_03525_));
 sky130_fd_sc_hd__nand2_1 _10505_ (.A(net175),
    .B(net156),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _10506_ (.A(net176),
    .B(net145),
    .Y(_03527_));
 sky130_fd_sc_hd__xor2_2 _10507_ (.A(_03526_),
    .B(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__xor2_2 _10508_ (.A(_02906_),
    .B(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__xor2_4 _10509_ (.A(_03525_),
    .B(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__a22oi_1 _10510_ (.A1(_00049_),
    .A2(_01562_),
    .B1(_02904_),
    .B2(_05115_),
    .Y(_03531_));
 sky130_fd_sc_hd__and4_2 _10511_ (.A(_05115_),
    .B(_00049_),
    .C(net197),
    .D(net198),
    .X(_03532_));
 sky130_fd_sc_hd__nor2_1 _10512_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__and4_1 _10513_ (.A(_00058_),
    .B(_00489_),
    .C(_00481_),
    .D(_01002_),
    .X(_03534_));
 sky130_fd_sc_hd__and4_1 _10514_ (.A(_00047_),
    .B(net196),
    .C(_02911_),
    .D(_02912_),
    .X(_03536_));
 sky130_fd_sc_hd__a22o_1 _10515_ (.A1(_00480_),
    .A2(net187),
    .B1(net188),
    .B2(_00989_),
    .X(_03537_));
 sky130_fd_sc_hd__nand4_2 _10516_ (.A(_00989_),
    .B(_00480_),
    .C(net187),
    .D(net188),
    .Y(_03538_));
 sky130_fd_sc_hd__and2_1 _10517_ (.A(net186),
    .B(net196),
    .X(_03539_));
 sky130_fd_sc_hd__a21o_1 _10518_ (.A1(_03537_),
    .A2(_03538_),
    .B1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__nand3_1 _10519_ (.A(_03537_),
    .B(_03538_),
    .C(_03539_),
    .Y(_03541_));
 sky130_fd_sc_hd__o211ai_2 _10520_ (.A1(_03534_),
    .A2(_03536_),
    .B1(_03540_),
    .C1(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__a211o_1 _10521_ (.A1(_03540_),
    .A2(_03541_),
    .B1(_03534_),
    .C1(_03536_),
    .X(_03543_));
 sky130_fd_sc_hd__nand3_1 _10522_ (.A(_03533_),
    .B(_03542_),
    .C(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21o_1 _10523_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03533_),
    .X(_03545_));
 sky130_fd_sc_hd__a21bo_1 _10524_ (.A1(_02907_),
    .A2(_02916_),
    .B1_N(_02915_),
    .X(_03547_));
 sky130_fd_sc_hd__and3_1 _10525_ (.A(_03544_),
    .B(_03545_),
    .C(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__a21o_1 _10526_ (.A1(_03544_),
    .A2(_03545_),
    .B1(_03547_),
    .X(_03549_));
 sky130_fd_sc_hd__and2b_1 _10527_ (.A_N(_03548_),
    .B(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__xor2_4 _10528_ (.A(_03530_),
    .B(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__and2_1 _10529_ (.A(_02931_),
    .B(_02935_),
    .X(_03552_));
 sky130_fd_sc_hd__a21o_1 _10530_ (.A1(_02930_),
    .A2(_02936_),
    .B1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a211oi_1 _10531_ (.A1(_02960_),
    .A2(_02961_),
    .B1(_02956_),
    .C1(_02277_),
    .Y(_03554_));
 sky130_fd_sc_hd__o21ai_2 _10532_ (.A1(_02955_),
    .A2(_03554_),
    .B1(_02962_),
    .Y(_03555_));
 sky130_fd_sc_hd__a22o_1 _10533_ (.A1(_01023_),
    .A2(_02950_),
    .B1(_02952_),
    .B2(_02953_),
    .X(_03556_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_03348_),
    .B(_01584_),
    .Y(_03558_));
 sky130_fd_sc_hd__and3_1 _10535_ (.A(net193),
    .B(_02239_),
    .C(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__xor2_2 _10536_ (.A(_03556_),
    .B(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__xor2_2 _10537_ (.A(_03555_),
    .B(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__xnor2_2 _10538_ (.A(_03553_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__nor2_1 _10539_ (.A(_02929_),
    .B(_02937_),
    .Y(_03563_));
 sky130_fd_sc_hd__a21oi_2 _10540_ (.A1(_02926_),
    .A2(_02938_),
    .B1(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xor2_2 _10541_ (.A(_03562_),
    .B(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__xor2_2 _10542_ (.A(_03551_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__xnor2_2 _10543_ (.A(_03523_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_4 _10544_ (.A(_03521_),
    .B(_03567_),
    .Y(_03569_));
 sky130_fd_sc_hd__and2b_1 _10545_ (.A_N(_02974_),
    .B(_02973_),
    .X(_03570_));
 sky130_fd_sc_hd__a21o_2 _10546_ (.A1(_02966_),
    .A2(_02975_),
    .B1(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__a21oi_4 _10547_ (.A1(_02980_),
    .A2(_03000_),
    .B1(_02999_),
    .Y(_03572_));
 sky130_fd_sc_hd__a22oi_1 _10548_ (.A1(_00507_),
    .A2(net231),
    .B1(_01603_),
    .B2(_00080_),
    .Y(_03573_));
 sky130_fd_sc_hd__and4_1 _10549_ (.A(net220),
    .B(net221),
    .C(net231),
    .D(net232),
    .X(_03574_));
 sky130_fd_sc_hd__nor2_2 _10550_ (.A(_03573_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_2 _10551_ (.A(_04752_),
    .B(net233),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_4 _10552_ (.A(_03575_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__a22o_1 _10553_ (.A1(net229),
    .A2(net224),
    .B1(net225),
    .B2(net228),
    .X(_03578_));
 sky130_fd_sc_hd__buf_2 _10554_ (.A(net225),
    .X(_03580_));
 sky130_fd_sc_hd__nand4_2 _10555_ (.A(_04741_),
    .B(_00086_),
    .C(net224),
    .D(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__and2_1 _10556_ (.A(net230),
    .B(net222),
    .X(_03582_));
 sky130_fd_sc_hd__a21o_1 _10557_ (.A1(_03578_),
    .A2(_03581_),
    .B1(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__nand3_1 _10558_ (.A(_03578_),
    .B(_03581_),
    .C(_03582_),
    .Y(_03584_));
 sky130_fd_sc_hd__a21bo_1 _10559_ (.A1(_02957_),
    .A2(_02959_),
    .B1_N(_02958_),
    .X(_03585_));
 sky130_fd_sc_hd__and3_1 _10560_ (.A(_03583_),
    .B(_03584_),
    .C(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__a21o_1 _10561_ (.A1(_03583_),
    .A2(_03584_),
    .B1(_03585_),
    .X(_03587_));
 sky130_fd_sc_hd__and2b_1 _10562_ (.A_N(_03586_),
    .B(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__xnor2_4 _10563_ (.A(_03577_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__o21bai_4 _10564_ (.A1(_02982_),
    .A2(_02985_),
    .B1_N(_02983_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand2_2 _10565_ (.A(_04906_),
    .B(net49),
    .Y(_03592_));
 sky130_fd_sc_hd__xnor2_4 _10566_ (.A(_03591_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__xnor2_4 _10567_ (.A(_02969_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__inv_2 _10568_ (.A(_02969_),
    .Y(_03595_));
 sky130_fd_sc_hd__a32o_2 _10569_ (.A1(_02968_),
    .A2(_03595_),
    .A3(_02970_),
    .B1(_02972_),
    .B2(_02967_),
    .X(_03596_));
 sky130_fd_sc_hd__xor2_4 _10570_ (.A(_03594_),
    .B(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__xnor2_4 _10571_ (.A(_03589_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__xor2_4 _10572_ (.A(_03572_),
    .B(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__xor2_4 _10573_ (.A(_03571_),
    .B(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__or2b_2 _10574_ (.A(_02994_),
    .B_N(_02996_),
    .X(_03602_));
 sky130_fd_sc_hd__and3_1 _10575_ (.A(_03004_),
    .B(_03005_),
    .C(_03007_),
    .X(_03603_));
 sky130_fd_sc_hd__a22oi_1 _10576_ (.A1(_00530_),
    .A2(_01068_),
    .B1(_01051_),
    .B2(_00543_),
    .Y(_03604_));
 sky130_fd_sc_hd__and4_1 _10577_ (.A(net37),
    .B(net46),
    .C(net38),
    .D(net47),
    .X(_03605_));
 sky130_fd_sc_hd__nor2_1 _10578_ (.A(_03604_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand2_1 _10579_ (.A(_00107_),
    .B(_01629_),
    .Y(_03607_));
 sky130_fd_sc_hd__xor2_1 _10580_ (.A(_03606_),
    .B(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__a22oi_1 _10581_ (.A1(_00097_),
    .A2(_01653_),
    .B1(_02329_),
    .B2(_04862_),
    .Y(_03609_));
 sky130_fd_sc_hd__and4_1 _10582_ (.A(_04862_),
    .B(net44),
    .C(net39),
    .D(net40),
    .X(_03610_));
 sky130_fd_sc_hd__nor2_1 _10583_ (.A(_03609_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21bo_1 _10584_ (.A1(_02988_),
    .A2(_02990_),
    .B1_N(_02989_),
    .X(_03613_));
 sky130_fd_sc_hd__xor2_1 _10585_ (.A(_03611_),
    .B(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__xnor2_1 _10586_ (.A(_03608_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__o21a_1 _10587_ (.A1(_03603_),
    .A2(_03011_),
    .B1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__or3_1 _10588_ (.A(_03603_),
    .B(_03011_),
    .C(_03615_),
    .X(_03617_));
 sky130_fd_sc_hd__or2b_2 _10589_ (.A(_03616_),
    .B_N(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__xnor2_4 _10590_ (.A(_03602_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__and4_1 _10591_ (.A(_03095_),
    .B(_04939_),
    .C(_01652_),
    .D(_03006_),
    .X(_03620_));
 sky130_fd_sc_hd__a32o_1 _10592_ (.A1(_00549_),
    .A2(net45),
    .A3(_03015_),
    .B1(_03014_),
    .B2(_01666_),
    .X(_03621_));
 sky130_fd_sc_hd__a22oi_1 _10593_ (.A1(_00549_),
    .A2(net56),
    .B1(net67),
    .B2(_04939_),
    .Y(_03622_));
 sky130_fd_sc_hd__and4_2 _10594_ (.A(_04939_),
    .B(_00549_),
    .C(net56),
    .D(net67),
    .X(_03624_));
 sky130_fd_sc_hd__nor2_1 _10595_ (.A(_03622_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__xor2_1 _10596_ (.A(_03621_),
    .B(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__nor2_1 _10597_ (.A(_03620_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__and2_1 _10598_ (.A(_03620_),
    .B(_03626_),
    .X(_03628_));
 sky130_fd_sc_hd__nor2_2 _10599_ (.A(_03627_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a22o_1 _10600_ (.A1(net34),
    .A2(net212),
    .B1(net223),
    .B2(_00109_),
    .X(_03630_));
 sky130_fd_sc_hd__nand4_1 _10601_ (.A(_00109_),
    .B(_00544_),
    .C(net212),
    .D(net223),
    .Y(_03631_));
 sky130_fd_sc_hd__and2_1 _10602_ (.A(_00550_),
    .B(net45),
    .X(_03632_));
 sky130_fd_sc_hd__a21o_1 _10603_ (.A1(_03630_),
    .A2(_03631_),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__nand3_1 _10604_ (.A(_03630_),
    .B(_03631_),
    .C(_03632_),
    .Y(_03635_));
 sky130_fd_sc_hd__nand2_1 _10605_ (.A(_03106_),
    .B(net223),
    .Y(_03636_));
 sky130_fd_sc_hd__and3_1 _10606_ (.A(net12),
    .B(net234),
    .C(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__a21oi_1 _10607_ (.A1(_03633_),
    .A2(_03635_),
    .B1(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__and3_1 _10608_ (.A(_03633_),
    .B(_03635_),
    .C(_03637_),
    .X(_03639_));
 sky130_fd_sc_hd__nor2_1 _10609_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__and2_1 _10610_ (.A(_03023_),
    .B(_03024_),
    .X(_03641_));
 sky130_fd_sc_hd__a21oi_2 _10611_ (.A1(_03018_),
    .A2(_03025_),
    .B1(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__xnor2_2 _10612_ (.A(_03640_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__xor2_4 _10613_ (.A(_03629_),
    .B(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(_03026_),
    .B(_03027_),
    .X(_03646_));
 sky130_fd_sc_hd__a21o_2 _10615_ (.A1(_03013_),
    .A2(_03028_),
    .B1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__xor2_4 _10616_ (.A(_03644_),
    .B(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__xor2_4 _10617_ (.A(_03619_),
    .B(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__and2_1 _10618_ (.A(_03029_),
    .B(_03030_),
    .X(_03650_));
 sky130_fd_sc_hd__a21oi_2 _10619_ (.A1(_03002_),
    .A2(_03032_),
    .B1(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__xnor2_4 _10620_ (.A(_03649_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_4 _10621_ (.A(_03600_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__and2b_1 _10622_ (.A_N(_03035_),
    .B(_03033_),
    .X(_03654_));
 sky130_fd_sc_hd__a21o_1 _10623_ (.A1(_02979_),
    .A2(_03036_),
    .B1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__xnor2_4 _10624_ (.A(_03653_),
    .B(_03655_),
    .Y(_03657_));
 sky130_fd_sc_hd__xnor2_4 _10625_ (.A(_03569_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__and2b_1 _10626_ (.A_N(_03039_),
    .B(_03037_),
    .X(_03659_));
 sky130_fd_sc_hd__a21oi_2 _10627_ (.A1(_02947_),
    .A2(_03040_),
    .B1(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__xor2_4 _10628_ (.A(_03658_),
    .B(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__xnor2_4 _10629_ (.A(_03519_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nor2_1 _10630_ (.A(_03041_),
    .B(_03043_),
    .Y(_03663_));
 sky130_fd_sc_hd__a21oi_2 _10631_ (.A1(_02890_),
    .A2(_03044_),
    .B1(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__xor2_4 _10632_ (.A(_03662_),
    .B(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__xnor2_4 _10633_ (.A(_03431_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__and2b_1 _10634_ (.A_N(_03045_),
    .B(_03046_),
    .X(_03668_));
 sky130_fd_sc_hd__a21oi_2 _10635_ (.A1(_02793_),
    .A2(_03047_),
    .B1(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__xor2_4 _10636_ (.A(_03666_),
    .B(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__xnor2_4 _10637_ (.A(_03316_),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__nor2_1 _10638_ (.A(_03048_),
    .B(_03049_),
    .Y(_03672_));
 sky130_fd_sc_hd__a21oi_4 _10639_ (.A1(_02666_),
    .A2(_03050_),
    .B1(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__xor2_2 _10640_ (.A(_03671_),
    .B(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__xnor2_2 _10641_ (.A(_03125_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nor2_1 _10642_ (.A(_03051_),
    .B(_03052_),
    .Y(_03676_));
 sky130_fd_sc_hd__a21oi_2 _10643_ (.A1(_02451_),
    .A2(_03054_),
    .B1(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__xor2_2 _10644_ (.A(_03675_),
    .B(_03677_),
    .X(_03679_));
 sky130_fd_sc_hd__xnor2_1 _10645_ (.A(_03079_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__a21oi_1 _10646_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__and3_1 _10647_ (.A(_03076_),
    .B(_03077_),
    .C(_03680_),
    .X(_03682_));
 sky130_fd_sc_hd__nor2_1 _10648_ (.A(_03681_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__xor2_1 _10649_ (.A(_03075_),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__nor2_1 _10650_ (.A(net285),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__and2_1 _10651_ (.A(net285),
    .B(_03684_),
    .X(_03686_));
 sky130_fd_sc_hd__nor2_1 _10652_ (.A(_03685_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__a21o_1 _10653_ (.A1(_03068_),
    .A2(_03071_),
    .B1(_03067_),
    .X(_03688_));
 sky130_fd_sc_hd__a21oi_1 _10654_ (.A1(_03687_),
    .A2(_03688_),
    .B1(_00166_),
    .Y(_03690_));
 sky130_fd_sc_hd__o21a_1 _10655_ (.A1(_03687_),
    .A2(_03688_),
    .B1(_03690_),
    .X(_00009_));
 sky130_fd_sc_hd__inv_2 _10656_ (.A(_03685_),
    .Y(_03691_));
 sky130_fd_sc_hd__a211o_1 _10657_ (.A1(_03070_),
    .A2(_03071_),
    .B1(_03686_),
    .C1(_03067_),
    .X(_03692_));
 sky130_fd_sc_hd__or2b_1 _10658_ (.A(_03123_),
    .B_N(_03082_),
    .X(_03693_));
 sky130_fd_sc_hd__or2b_1 _10659_ (.A(_03124_),
    .B_N(_03081_),
    .X(_03694_));
 sky130_fd_sc_hd__nand2_2 _10660_ (.A(_03693_),
    .B(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__or2b_1 _10661_ (.A(_03089_),
    .B_N(_03121_),
    .X(_03696_));
 sky130_fd_sc_hd__a21bo_2 _10662_ (.A1(_03086_),
    .A2(_03122_),
    .B1_N(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__and2b_1 _10663_ (.A_N(_03313_),
    .B(_03129_),
    .X(_03698_));
 sky130_fd_sc_hd__a21o_2 _10664_ (.A1(_03126_),
    .A2(_03314_),
    .B1(_03698_),
    .X(_03700_));
 sky130_fd_sc_hd__and2b_1 _10665_ (.A_N(_03090_),
    .B(_03120_),
    .X(_03701_));
 sky130_fd_sc_hd__or2_2 _10666_ (.A(_03118_),
    .B(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__o21ba_2 _10667_ (.A1(_03158_),
    .A2(_03246_),
    .B1_N(_03245_),
    .X(_03703_));
 sky130_fd_sc_hd__o21ba_2 _10668_ (.A1(_03113_),
    .A2(_03115_),
    .B1_N(_03112_),
    .X(_03704_));
 sky130_fd_sc_hd__or2b_1 _10669_ (.A(_03132_),
    .B_N(_03156_),
    .X(_03705_));
 sky130_fd_sc_hd__or2b_1 _10670_ (.A(_03157_),
    .B_N(_03131_),
    .X(_03706_));
 sky130_fd_sc_hd__and2_1 _10671_ (.A(_02466_),
    .B(_03100_),
    .X(_03707_));
 sky130_fd_sc_hd__and2b_1 _10672_ (.A_N(_03101_),
    .B(_03102_),
    .X(_03708_));
 sky130_fd_sc_hd__and2_1 _10673_ (.A(net170),
    .B(_01188_),
    .X(_03709_));
 sky130_fd_sc_hd__a21oi_1 _10674_ (.A1(_06227_),
    .A2(_02464_),
    .B1(_03709_),
    .Y(_03711_));
 sky130_fd_sc_hd__and3_1 _10675_ (.A(_06227_),
    .B(net164),
    .C(_03709_),
    .X(_03712_));
 sky130_fd_sc_hd__o2bb2a_1 _10676_ (.A1_N(_01777_),
    .A2_N(_00617_),
    .B1(_03711_),
    .B2(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__and4bb_1 _10677_ (.A_N(_03711_),
    .B_N(_03712_),
    .C(_01777_),
    .D(_00617_),
    .X(_03714_));
 sky130_fd_sc_hd__or2_1 _10678_ (.A(_03713_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__o21a_1 _10679_ (.A1(_03098_),
    .A2(_03099_),
    .B1(_03097_),
    .X(_03716_));
 sky130_fd_sc_hd__or2_1 _10680_ (.A(_03715_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_03715_),
    .B(_03716_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _10682_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__o21bai_1 _10683_ (.A1(_03707_),
    .A2(_03708_),
    .B1_N(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__or3b_1 _10684_ (.A(_03707_),
    .B(_03708_),
    .C_N(_03719_),
    .X(_03722_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(_03720_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_00270_),
    .B(_01157_),
    .Y(_03724_));
 sky130_fd_sc_hd__xor2_1 _10687_ (.A(_03723_),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__o21a_1 _10688_ (.A1(_03104_),
    .A2(_03110_),
    .B1(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nor3_1 _10689_ (.A(_03104_),
    .B(_03110_),
    .C(_03725_),
    .Y(_03727_));
 sky130_fd_sc_hd__nor2_1 _10690_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand2_1 _10691_ (.A(_06243_),
    .B(net173),
    .Y(_03729_));
 sky130_fd_sc_hd__xor2_1 _10692_ (.A(_03728_),
    .B(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__a21oi_1 _10693_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__and3_1 _10694_ (.A(_03705_),
    .B(_03706_),
    .C(_03730_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_2 _10695_ (.A(_03731_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_4 _10696_ (.A(_03704_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__xnor2_4 _10697_ (.A(_03703_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__xnor2_4 _10698_ (.A(_03702_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__xor2_2 _10699_ (.A(_03700_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__xnor2_2 _10700_ (.A(_03697_),
    .B(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__a21o_2 _10701_ (.A1(_03248_),
    .A2(_03312_),
    .B1(_03310_),
    .X(_03740_));
 sky130_fd_sc_hd__a21o_1 _10702_ (.A1(_03317_),
    .A2(_03430_),
    .B1(_03428_),
    .X(_03741_));
 sky130_fd_sc_hd__and2b_1 _10703_ (.A_N(_03154_),
    .B(_03136_),
    .X(_03742_));
 sky130_fd_sc_hd__a21oi_4 _10704_ (.A1(_03135_),
    .A2(_03155_),
    .B1(_03742_),
    .Y(_03744_));
 sky130_fd_sc_hd__or2b_1 _10705_ (.A(_03187_),
    .B_N(_03202_),
    .X(_03745_));
 sky130_fd_sc_hd__o21a_2 _10706_ (.A1(_03200_),
    .A2(_03201_),
    .B1(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__a21oi_2 _10707_ (.A1(_03138_),
    .A2(_03153_),
    .B1(_03151_),
    .Y(_03747_));
 sky130_fd_sc_hd__a21oi_2 _10708_ (.A1(_03170_),
    .A2(_03186_),
    .B1(_03184_),
    .Y(_03748_));
 sky130_fd_sc_hd__and2b_1 _10709_ (.A_N(_03146_),
    .B(_03147_),
    .X(_03749_));
 sky130_fd_sc_hd__a31oi_2 _10710_ (.A1(_06130_),
    .A2(_02464_),
    .A3(_03148_),
    .B1(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__a21o_1 _10711_ (.A1(_02500_),
    .A2(_03166_),
    .B1(_03168_),
    .X(_03751_));
 sky130_fd_sc_hd__a22o_1 _10712_ (.A1(net20),
    .A2(net29),
    .B1(net30),
    .B2(net19),
    .X(_03752_));
 sky130_fd_sc_hd__nand4_1 _10713_ (.A(net19),
    .B(_00706_),
    .C(_00647_),
    .D(_01181_),
    .Y(_03753_));
 sky130_fd_sc_hd__a22oi_2 _10714_ (.A1(_06261_),
    .A2(_01784_),
    .B1(_03752_),
    .B2(_03753_),
    .Y(_03755_));
 sky130_fd_sc_hd__and4_1 _10715_ (.A(_06261_),
    .B(net31),
    .C(_03752_),
    .D(_03753_),
    .X(_03756_));
 sky130_fd_sc_hd__o21ai_1 _10716_ (.A1(_03144_),
    .A2(_03145_),
    .B1(_03143_),
    .Y(_03757_));
 sky130_fd_sc_hd__or3b_1 _10717_ (.A(_03755_),
    .B(_03756_),
    .C_N(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10718_ (.A(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__o21bai_2 _10719_ (.A1(_03755_),
    .A2(_03756_),
    .B1_N(_03757_),
    .Y(_03760_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_03759_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__xnor2_1 _10721_ (.A(_03751_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_1 _10722_ (.A(_03750_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__xnor2_2 _10723_ (.A(_03748_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__xnor2_2 _10724_ (.A(_03747_),
    .B(_03764_),
    .Y(_03766_));
 sky130_fd_sc_hd__xnor2_4 _10725_ (.A(_03746_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__xnor2_4 _10726_ (.A(_03744_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nor2_1 _10727_ (.A(_03237_),
    .B(_03240_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand3_1 _10728_ (.A(_00250_),
    .B(_00706_),
    .C(_03164_),
    .Y(_03770_));
 sky130_fd_sc_hd__a22oi_1 _10729_ (.A1(_00250_),
    .A2(_01217_),
    .B1(_02498_),
    .B2(_06264_),
    .Y(_03771_));
 sky130_fd_sc_hd__and4_1 _10730_ (.A(_06264_),
    .B(_00250_),
    .C(_01217_),
    .D(_02498_),
    .X(_03772_));
 sky130_fd_sc_hd__or2_1 _10731_ (.A(_03771_),
    .B(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__a21o_1 _10732_ (.A1(_03163_),
    .A2(_03770_),
    .B1(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__nand3_1 _10733_ (.A(_03163_),
    .B(_03770_),
    .C(_03773_),
    .Y(_03775_));
 sky130_fd_sc_hd__and2_1 _10734_ (.A(_03774_),
    .B(_03775_),
    .X(_03777_));
 sky130_fd_sc_hd__and2b_1 _10735_ (.A_N(_03177_),
    .B(_03178_),
    .X(_03778_));
 sky130_fd_sc_hd__and3_1 _10736_ (.A(_06159_),
    .B(_03180_),
    .C(_03179_),
    .X(_03779_));
 sky130_fd_sc_hd__a22oi_2 _10737_ (.A1(net91),
    .A2(_00703_),
    .B1(net92),
    .B2(_00238_),
    .Y(_03780_));
 sky130_fd_sc_hd__and4_1 _10738_ (.A(net98),
    .B(net91),
    .C(net99),
    .D(net92),
    .X(_03781_));
 sky130_fd_sc_hd__nor2_1 _10739_ (.A(_03780_),
    .B(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _10740_ (.A(_00200_),
    .B(net101),
    .Y(_03783_));
 sky130_fd_sc_hd__xnor2_1 _10741_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__o21a_1 _10742_ (.A1(_03174_),
    .A2(_03176_),
    .B1(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__nor3_1 _10743_ (.A(_03174_),
    .B(_03176_),
    .C(_03784_),
    .Y(_03786_));
 sky130_fd_sc_hd__nor2_1 _10744_ (.A(_03785_),
    .B(_03786_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_06284_),
    .B(net102),
    .Y(_03789_));
 sky130_fd_sc_hd__xnor2_1 _10746_ (.A(_03788_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__o21a_1 _10747_ (.A1(_03778_),
    .A2(_03779_),
    .B1(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__or3_1 _10748_ (.A(_03778_),
    .B(_03779_),
    .C(_03790_),
    .X(_03792_));
 sky130_fd_sc_hd__and2b_1 _10749_ (.A_N(_03791_),
    .B(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__xor2_2 _10750_ (.A(_03777_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__and2_1 _10751_ (.A(_02546_),
    .B(_03193_),
    .X(_03795_));
 sky130_fd_sc_hd__a21o_1 _10752_ (.A1(_03190_),
    .A2(_03195_),
    .B1(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__a21boi_2 _10753_ (.A1(_03213_),
    .A2(_03223_),
    .B1_N(_03222_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _10754_ (.A(_06253_),
    .B(_01858_),
    .Y(_03799_));
 sky130_fd_sc_hd__a21oi_1 _10755_ (.A1(_06134_),
    .A2(_01251_),
    .B1(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__xnor2_1 _10756_ (.A(_03212_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__xor2_1 _10757_ (.A(_03797_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__nand2_1 _10758_ (.A(_03796_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__or2_1 _10759_ (.A(_03796_),
    .B(_03802_),
    .X(_03804_));
 sky130_fd_sc_hd__nand2_1 _10760_ (.A(_03803_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__a21oi_1 _10761_ (.A1(_03188_),
    .A2(_03198_),
    .B1(_03197_),
    .Y(_03806_));
 sky130_fd_sc_hd__nor2_1 _10762_ (.A(_03805_),
    .B(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__and2_1 _10763_ (.A(_03805_),
    .B(_03806_),
    .X(_03808_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(_03807_),
    .B(_03808_),
    .Y(_03810_));
 sky130_fd_sc_hd__xnor2_1 _10765_ (.A(_03794_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__nor2_1 _10766_ (.A(_03228_),
    .B(_03233_),
    .Y(_03812_));
 sky130_fd_sc_hd__nand2_1 _10767_ (.A(_03228_),
    .B(_03233_),
    .Y(_03813_));
 sky130_fd_sc_hd__o21ai_1 _10768_ (.A1(_03225_),
    .A2(_03812_),
    .B1(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__a21o_1 _10769_ (.A1(_03255_),
    .A2(_03275_),
    .B1(_03274_),
    .X(_03815_));
 sky130_fd_sc_hd__a22oi_2 _10770_ (.A1(_00210_),
    .A2(_01250_),
    .B1(_03210_),
    .B2(_06274_),
    .Y(_03816_));
 sky130_fd_sc_hd__and4_1 _10771_ (.A(_06274_),
    .B(_00210_),
    .C(_01250_),
    .D(net138),
    .X(_03817_));
 sky130_fd_sc_hd__or2_1 _10772_ (.A(_03816_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__a22o_1 _10773_ (.A1(net135),
    .A2(net128),
    .B1(net129),
    .B2(net133),
    .X(_03819_));
 sky130_fd_sc_hd__nand4_1 _10774_ (.A(net133),
    .B(net135),
    .C(net128),
    .D(net129),
    .Y(_03821_));
 sky130_fd_sc_hd__and2_1 _10775_ (.A(net127),
    .B(net136),
    .X(_03822_));
 sky130_fd_sc_hd__a21o_1 _10776_ (.A1(_03819_),
    .A2(_03821_),
    .B1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__nand3_1 _10777_ (.A(_03819_),
    .B(_03821_),
    .C(_03822_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21bo_1 _10778_ (.A1(_03217_),
    .A2(_03219_),
    .B1_N(_03218_),
    .X(_03825_));
 sky130_fd_sc_hd__and3_1 _10779_ (.A(_03823_),
    .B(_03824_),
    .C(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__a21oi_1 _10780_ (.A1(_03823_),
    .A2(_03824_),
    .B1(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__or2_2 _10781_ (.A(_03826_),
    .B(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__xnor2_2 _10782_ (.A(_03818_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__a32o_1 _10783_ (.A1(_06178_),
    .A2(_02592_),
    .A3(_03258_),
    .B1(_03257_),
    .B2(_00749_),
    .X(_03830_));
 sky130_fd_sc_hd__or2b_1 _10784_ (.A(_03230_),
    .B_N(_03231_),
    .X(_03832_));
 sky130_fd_sc_hd__and3_1 _10785_ (.A(_06151_),
    .B(_01872_),
    .C(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__xnor2_2 _10786_ (.A(_03830_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__xor2_1 _10787_ (.A(_03829_),
    .B(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__xor2_1 _10788_ (.A(_03815_),
    .B(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__xnor2_1 _10789_ (.A(_03814_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__and2b_1 _10790_ (.A_N(_03209_),
    .B(_03235_),
    .X(_03838_));
 sky130_fd_sc_hd__a21oi_1 _10791_ (.A1(_03207_),
    .A2(_03236_),
    .B1(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__or2_1 _10792_ (.A(_03837_),
    .B(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__nand2_1 _10793_ (.A(_03837_),
    .B(_03839_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_03840_),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__xor2_1 _10795_ (.A(_03811_),
    .B(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__o21a_1 _10796_ (.A1(_03769_),
    .A2(_03242_),
    .B1(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__nor3_1 _10797_ (.A(_03769_),
    .B(_03242_),
    .C(_03844_),
    .Y(_03846_));
 sky130_fd_sc_hd__nor2_2 _10798_ (.A(_03845_),
    .B(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__xor2_4 _10799_ (.A(_03768_),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__and2b_1 _10800_ (.A_N(_03305_),
    .B(_03253_),
    .X(_03849_));
 sky130_fd_sc_hd__a21o_1 _10801_ (.A1(_03254_),
    .A2(_03303_),
    .B1(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__or2_1 _10802_ (.A(_03380_),
    .B(_03383_),
    .X(_03851_));
 sky130_fd_sc_hd__o21ai_2 _10803_ (.A1(_03335_),
    .A2(_03384_),
    .B1(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__and2b_1 _10804_ (.A_N(_03301_),
    .B(_03300_),
    .X(_03854_));
 sky130_fd_sc_hd__a21o_1 _10805_ (.A1(_03277_),
    .A2(_03302_),
    .B1(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__and2b_1 _10806_ (.A_N(_03333_),
    .B(_03321_),
    .X(_03856_));
 sky130_fd_sc_hd__a21o_1 _10807_ (.A1(_03320_),
    .A2(_03334_),
    .B1(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(_03269_),
    .B(_03272_),
    .Y(_03858_));
 sky130_fd_sc_hd__clkbuf_4 _10809_ (.A(net216),
    .X(_03859_));
 sky130_fd_sc_hd__and3_1 _10810_ (.A(_06086_),
    .B(_03859_),
    .C(_03279_),
    .X(_03860_));
 sky130_fd_sc_hd__and3_1 _10811_ (.A(net143),
    .B(net144),
    .C(net154),
    .X(_03861_));
 sky130_fd_sc_hd__a22o_1 _10812_ (.A1(net144),
    .A2(net153),
    .B1(net154),
    .B2(net143),
    .X(_03862_));
 sky130_fd_sc_hd__a21bo_1 _10813_ (.A1(net153),
    .A2(_03861_),
    .B1_N(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_06311_),
    .B(net155),
    .Y(_03865_));
 sky130_fd_sc_hd__xor2_1 _10815_ (.A(_03863_),
    .B(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__a22o_1 _10816_ (.A1(_01293_),
    .A2(net146),
    .B1(_02615_),
    .B2(_06319_),
    .X(_03867_));
 sky130_fd_sc_hd__nand4_2 _10817_ (.A(_06319_),
    .B(_01293_),
    .C(_01309_),
    .D(_02615_),
    .Y(_03868_));
 sky130_fd_sc_hd__nand2_1 _10818_ (.A(_03867_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__a21bo_1 _10819_ (.A1(_03263_),
    .A2(_03265_),
    .B1_N(_03264_),
    .X(_03870_));
 sky130_fd_sc_hd__xnor2_1 _10820_ (.A(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__xor2_1 _10821_ (.A(_03866_),
    .B(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__o21ai_1 _10822_ (.A1(_03860_),
    .A2(_03284_),
    .B1(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__or3_1 _10823_ (.A(_03860_),
    .B(_03284_),
    .C(_03872_),
    .X(_03874_));
 sky130_fd_sc_hd__and3_1 _10824_ (.A(_03858_),
    .B(_03873_),
    .C(_03874_),
    .X(_03876_));
 sky130_fd_sc_hd__a21oi_1 _10825_ (.A1(_03873_),
    .A2(_03874_),
    .B1(_03858_),
    .Y(_03877_));
 sky130_fd_sc_hd__nor2_2 _10826_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__and3_1 _10827_ (.A(_06362_),
    .B(_02626_),
    .C(_03288_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _10828_ (.A(_06362_),
    .B(_03859_),
    .Y(_03880_));
 sky130_fd_sc_hd__o21ba_1 _10829_ (.A1(_03287_),
    .A2(_03879_),
    .B1_N(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__nor3b_1 _10830_ (.A(_03287_),
    .B(_03879_),
    .C_N(_03880_),
    .Y(_03882_));
 sky130_fd_sc_hd__nor2_1 _10831_ (.A(_03881_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__a22o_1 _10832_ (.A1(_00810_),
    .A2(net214),
    .B1(net206),
    .B2(_00297_),
    .X(_03884_));
 sky130_fd_sc_hd__nand4_1 _10833_ (.A(_00297_),
    .B(_00810_),
    .C(_00757_),
    .D(_01365_),
    .Y(_03885_));
 sky130_fd_sc_hd__a22o_1 _10834_ (.A1(_00343_),
    .A2(net215),
    .B1(_03884_),
    .B2(_03885_),
    .X(_03887_));
 sky130_fd_sc_hd__nand4_1 _10835_ (.A(_00343_),
    .B(_02626_),
    .C(_03884_),
    .D(_03885_),
    .Y(_03888_));
 sky130_fd_sc_hd__nand2_1 _10836_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _10837_ (.A(_06173_),
    .B(_01365_),
    .Y(_03890_));
 sky130_fd_sc_hd__and3_1 _10838_ (.A(_06304_),
    .B(_01986_),
    .C(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__xor2_2 _10839_ (.A(_03889_),
    .B(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _10840_ (.A(_03294_),
    .B(_03295_),
    .X(_03893_));
 sky130_fd_sc_hd__a21oi_2 _10841_ (.A1(_03290_),
    .A2(_03296_),
    .B1(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__xor2_2 _10842_ (.A(_03892_),
    .B(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__xor2_2 _10843_ (.A(_03883_),
    .B(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__nor2_1 _10844_ (.A(_03297_),
    .B(_03298_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _10845_ (.A(_03297_),
    .B(_03298_),
    .Y(_03899_));
 sky130_fd_sc_hd__o21a_1 _10846_ (.A1(_03285_),
    .A2(_03898_),
    .B1(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__xnor2_2 _10847_ (.A(_03896_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__xor2_2 _10848_ (.A(_03878_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__xnor2_2 _10849_ (.A(_03857_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__xnor2_2 _10850_ (.A(_03855_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__xor2_2 _10851_ (.A(_03852_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__xnor2_2 _10852_ (.A(_03850_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__or2b_1 _10853_ (.A(_03252_),
    .B_N(_03306_),
    .X(_03907_));
 sky130_fd_sc_hd__a21boi_2 _10854_ (.A1(_03250_),
    .A2(_03307_),
    .B1_N(_03907_),
    .Y(_03909_));
 sky130_fd_sc_hd__nor2_1 _10855_ (.A(_03906_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__and2_1 _10856_ (.A(_03906_),
    .B(_03909_),
    .X(_03911_));
 sky130_fd_sc_hd__nor2_1 _10857_ (.A(_03910_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__xnor2_2 _10858_ (.A(_03848_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__xnor2_2 _10859_ (.A(_03741_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__xor2_4 _10860_ (.A(_03740_),
    .B(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__or2b_1 _10861_ (.A(_03385_),
    .B_N(_03426_),
    .X(_03916_));
 sky130_fd_sc_hd__o21ai_4 _10862_ (.A1(_03422_),
    .A2(_03424_),
    .B1(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21boi_2 _10863_ (.A1(_03432_),
    .A2(_03516_),
    .B1_N(_03515_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor2_1 _10864_ (.A(_03324_),
    .B(_03331_),
    .Y(_03920_));
 sky130_fd_sc_hd__a21o_2 _10865_ (.A1(_03323_),
    .A2(_03332_),
    .B1(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__a21o_2 _10866_ (.A1(_03345_),
    .A2(_03360_),
    .B1(_03358_),
    .X(_03922_));
 sky130_fd_sc_hd__nor2_1 _10867_ (.A(_03325_),
    .B(_03329_),
    .Y(_03923_));
 sky130_fd_sc_hd__a21o_2 _10868_ (.A1(_02676_),
    .A2(_03330_),
    .B1(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__a31o_2 _10869_ (.A1(_03340_),
    .A2(_03341_),
    .A3(_03344_),
    .B1(_02697_),
    .X(_03925_));
 sky130_fd_sc_hd__a21bo_2 _10870_ (.A1(_03336_),
    .A2(_03339_),
    .B1_N(_03338_),
    .X(_03926_));
 sky130_fd_sc_hd__a22oi_1 _10871_ (.A1(_00834_),
    .A2(_01367_),
    .B1(_01987_),
    .B2(_06384_),
    .Y(_03927_));
 sky130_fd_sc_hd__and4_1 _10872_ (.A(net238),
    .B(_00834_),
    .C(net250),
    .D(net251),
    .X(_03928_));
 sky130_fd_sc_hd__nor2_2 _10873_ (.A(_03927_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__xnor2_4 _10874_ (.A(_03926_),
    .B(_03929_),
    .Y(_03931_));
 sky130_fd_sc_hd__xor2_4 _10875_ (.A(_03328_),
    .B(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__xnor2_4 _10876_ (.A(_03925_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__xnor2_4 _10877_ (.A(_03924_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__xor2_4 _10878_ (.A(_03922_),
    .B(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__xor2_4 _10879_ (.A(_03921_),
    .B(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__a22o_1 _10880_ (.A1(_00366_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_06383_),
    .X(_03937_));
 sky130_fd_sc_hd__and4_1 _10881_ (.A(_06383_),
    .B(_00366_),
    .C(_02694_),
    .D(net242),
    .X(_03938_));
 sky130_fd_sc_hd__inv_2 _10882_ (.A(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a22oi_1 _10883_ (.A1(_01385_),
    .A2(_00830_),
    .B1(_03937_),
    .B2(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__and4b_1 _10884_ (.A_N(_03938_),
    .B(_00830_),
    .C(_01385_),
    .D(_03937_),
    .X(_03942_));
 sky130_fd_sc_hd__or2_2 _10885_ (.A(_03940_),
    .B(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__a21bo_1 _10886_ (.A1(_03347_),
    .A2(_03350_),
    .B1_N(_03349_),
    .X(_03944_));
 sky130_fd_sc_hd__inv_2 _10887_ (.A(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__o21bai_1 _10888_ (.A1(_03366_),
    .A2(_03369_),
    .B1_N(_03367_),
    .Y(_03946_));
 sky130_fd_sc_hd__a22o_1 _10889_ (.A1(net3),
    .A2(net11),
    .B1(net13),
    .B2(net2),
    .X(_03947_));
 sky130_fd_sc_hd__nand4_2 _10890_ (.A(_00357_),
    .B(net3),
    .C(net11),
    .D(net13),
    .Y(_03948_));
 sky130_fd_sc_hd__a22o_1 _10891_ (.A1(_06375_),
    .A2(net14),
    .B1(_03947_),
    .B2(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand4_2 _10892_ (.A(_06375_),
    .B(_02019_),
    .C(_03947_),
    .D(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__and3_1 _10893_ (.A(_03946_),
    .B(_03949_),
    .C(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__a21oi_1 _10894_ (.A1(_03949_),
    .A2(_03950_),
    .B1(_03946_),
    .Y(_03953_));
 sky130_fd_sc_hd__or3_1 _10895_ (.A(_03945_),
    .B(_03951_),
    .C(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__o21ai_1 _10896_ (.A1(_03951_),
    .A2(_03953_),
    .B1(_03945_),
    .Y(_03955_));
 sky130_fd_sc_hd__a21bo_1 _10897_ (.A1(_03346_),
    .A2(_03354_),
    .B1_N(_03353_),
    .X(_03956_));
 sky130_fd_sc_hd__and3_1 _10898_ (.A(_03954_),
    .B(_03955_),
    .C(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__a21oi_1 _10899_ (.A1(_03954_),
    .A2(_03955_),
    .B1(_03956_),
    .Y(_03958_));
 sky130_fd_sc_hd__nor2_1 _10900_ (.A(_03957_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__xnor2_2 _10901_ (.A(_03943_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__a22o_1 _10902_ (.A1(_05750_),
    .A2(_02733_),
    .B1(_03371_),
    .B2(_03372_),
    .X(_03961_));
 sky130_fd_sc_hd__a21oi_2 _10903_ (.A1(_03394_),
    .A2(_03401_),
    .B1(_03400_),
    .Y(_03962_));
 sky130_fd_sc_hd__a22o_1 _10904_ (.A1(_00822_),
    .A2(_01410_),
    .B1(_02731_),
    .B2(_06368_),
    .X(_03964_));
 sky130_fd_sc_hd__nand4_2 _10905_ (.A(_06368_),
    .B(_00822_),
    .C(_01410_),
    .D(_02731_),
    .Y(_03965_));
 sky130_fd_sc_hd__and4_2 _10906_ (.A(_06343_),
    .B(net66),
    .C(_03964_),
    .D(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__buf_2 _10907_ (.A(net66),
    .X(_03967_));
 sky130_fd_sc_hd__a22oi_1 _10908_ (.A1(_06343_),
    .A2(_03967_),
    .B1(_03964_),
    .B2(_03965_),
    .Y(_03968_));
 sky130_fd_sc_hd__or2_1 _10909_ (.A(_03966_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__xnor2_1 _10910_ (.A(_03962_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__xnor2_2 _10911_ (.A(_03961_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__and2_1 _10912_ (.A(_03365_),
    .B(_03374_),
    .X(_03972_));
 sky130_fd_sc_hd__a21oi_2 _10913_ (.A1(_03364_),
    .A2(_03375_),
    .B1(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_2 _10914_ (.A(_03971_),
    .B(_03973_),
    .Y(_03975_));
 sky130_fd_sc_hd__xor2_2 _10915_ (.A(_03960_),
    .B(_03975_),
    .X(_03976_));
 sky130_fd_sc_hd__nand2_1 _10916_ (.A(_03376_),
    .B(_03378_),
    .Y(_03977_));
 sky130_fd_sc_hd__a21boi_2 _10917_ (.A1(_03362_),
    .A2(_03379_),
    .B1_N(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__xnor2_2 _10918_ (.A(_03976_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__xor2_2 _10919_ (.A(_03936_),
    .B(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__and2b_1 _10920_ (.A_N(_03419_),
    .B(_03391_),
    .X(_03981_));
 sky130_fd_sc_hd__a21o_1 _10921_ (.A1(_03393_),
    .A2(_03418_),
    .B1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a21bo_1 _10922_ (.A1(_03450_),
    .A2(_03482_),
    .B1_N(_03481_),
    .X(_03983_));
 sky130_fd_sc_hd__or2_1 _10923_ (.A(_03412_),
    .B(_03416_),
    .X(_03984_));
 sky130_fd_sc_hd__o21ai_2 _10924_ (.A1(_03404_),
    .A2(_03417_),
    .B1(_03984_),
    .Y(_03986_));
 sky130_fd_sc_hd__a21oi_2 _10925_ (.A1(_03434_),
    .A2(_03448_),
    .B1(_03446_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_2 _10926_ (.A(_03397_),
    .B(_03399_),
    .Y(_03988_));
 sky130_fd_sc_hd__a22o_1 _10927_ (.A1(net55),
    .A2(net64),
    .B1(net57),
    .B2(net63),
    .X(_03989_));
 sky130_fd_sc_hd__nand4_2 _10928_ (.A(net63),
    .B(net55),
    .C(net64),
    .D(net57),
    .Y(_03990_));
 sky130_fd_sc_hd__a22o_1 _10929_ (.A1(_00387_),
    .A2(net65),
    .B1(_03989_),
    .B2(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__nand4_1 _10930_ (.A(_00387_),
    .B(net65),
    .C(_03989_),
    .D(_03990_),
    .Y(_03992_));
 sky130_fd_sc_hd__and3_1 _10931_ (.A(_03406_),
    .B(_03991_),
    .C(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__a21o_1 _10932_ (.A1(_03991_),
    .A2(_03992_),
    .B1(_03406_),
    .X(_03994_));
 sky130_fd_sc_hd__or2b_1 _10933_ (.A(_03993_),
    .B_N(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__xnor2_2 _10934_ (.A(_03988_),
    .B(_03995_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_2 _10935_ (.A(_06347_),
    .B(_02765_),
    .Y(_03998_));
 sky130_fd_sc_hd__and4_1 _10936_ (.A(net71),
    .B(net72),
    .C(net83),
    .D(net84),
    .X(_03999_));
 sky130_fd_sc_hd__and2_1 _10937_ (.A(_03409_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__a22oi_1 _10938_ (.A1(_00431_),
    .A2(_01443_),
    .B1(_02064_),
    .B2(_06424_),
    .Y(_04001_));
 sky130_fd_sc_hd__nor2_1 _10939_ (.A(_03409_),
    .B(_03999_),
    .Y(_04002_));
 sky130_fd_sc_hd__or3_2 _10940_ (.A(_04000_),
    .B(_04001_),
    .C(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__xor2_2 _10941_ (.A(_03998_),
    .B(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__and2_1 _10942_ (.A(_02773_),
    .B(_03409_),
    .X(_04005_));
 sky130_fd_sc_hd__a31o_1 _10943_ (.A1(_03407_),
    .A2(_03408_),
    .A3(_03410_),
    .B1(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__xor2_2 _10944_ (.A(_04004_),
    .B(_04006_),
    .X(_04008_));
 sky130_fd_sc_hd__xor2_2 _10945_ (.A(_03997_),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__xnor2_2 _10946_ (.A(_03987_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__xnor2_2 _10947_ (.A(_03986_),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__xnor2_2 _10948_ (.A(_03983_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__xnor2_2 _10949_ (.A(_03982_),
    .B(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__and2b_1 _10950_ (.A_N(_03388_),
    .B(_03420_),
    .X(_04014_));
 sky130_fd_sc_hd__a21oi_1 _10951_ (.A1(_03387_),
    .A2(_03421_),
    .B1(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__xor2_1 _10952_ (.A(_04013_),
    .B(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__xnor2_1 _10953_ (.A(_03980_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__nor2_1 _10954_ (.A(_03918_),
    .B(_04017_),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2_1 _10955_ (.A(_03918_),
    .B(_04017_),
    .Y(_04020_));
 sky130_fd_sc_hd__and2b_1 _10956_ (.A_N(_04019_),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__xor2_4 _10957_ (.A(_03917_),
    .B(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__or2b_2 _10958_ (.A(_03510_),
    .B_N(_03512_),
    .X(_04023_));
 sky130_fd_sc_hd__and2_1 _10959_ (.A(_03523_),
    .B(_03566_),
    .X(_04024_));
 sky130_fd_sc_hd__and2b_1 _10960_ (.A_N(_03567_),
    .B(_03521_),
    .X(_04025_));
 sky130_fd_sc_hd__nand2_2 _10961_ (.A(_03442_),
    .B(_03444_),
    .Y(_04026_));
 sky130_fd_sc_hd__o21ba_2 _10962_ (.A1(_03466_),
    .A2(_03474_),
    .B1_N(_03473_),
    .X(_04027_));
 sky130_fd_sc_hd__and3_1 _10963_ (.A(net80),
    .B(net81),
    .C(net74),
    .X(_04028_));
 sky130_fd_sc_hd__a22o_1 _10964_ (.A1(net81),
    .A2(net74),
    .B1(net75),
    .B2(net80),
    .X(_04030_));
 sky130_fd_sc_hd__a21bo_1 _10965_ (.A1(net75),
    .A2(_04028_),
    .B1_N(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__nand2_2 _10966_ (.A(_01487_),
    .B(_00937_),
    .Y(_04032_));
 sky130_fd_sc_hd__xor2_4 _10967_ (.A(_04031_),
    .B(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__and2_2 _10968_ (.A(_03439_),
    .B(_03441_),
    .X(_04034_));
 sky130_fd_sc_hd__xor2_4 _10969_ (.A(_04033_),
    .B(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__xor2_4 _10970_ (.A(_04027_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__xor2_4 _10971_ (.A(_04026_),
    .B(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__a22o_1 _10972_ (.A1(_00956_),
    .A2(_00910_),
    .B1(net119),
    .B2(_00454_),
    .X(_04038_));
 sky130_fd_sc_hd__nand4_1 _10973_ (.A(_00454_),
    .B(_00956_),
    .C(_00910_),
    .D(_01484_),
    .Y(_04039_));
 sky130_fd_sc_hd__and2_1 _10974_ (.A(_06437_),
    .B(_02132_),
    .X(_04041_));
 sky130_fd_sc_hd__a21oi_1 _10975_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__and3_1 _10976_ (.A(_04038_),
    .B(_04039_),
    .C(_04041_),
    .X(_04043_));
 sky130_fd_sc_hd__or2_2 _10977_ (.A(_04042_),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__a21boi_4 _10978_ (.A1(_03467_),
    .A2(_03470_),
    .B1_N(_03468_),
    .Y(_04045_));
 sky130_fd_sc_hd__xor2_4 _10979_ (.A(_04044_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__a22oi_2 _10980_ (.A1(_00438_),
    .A2(_01520_),
    .B1(_02164_),
    .B2(_06416_),
    .Y(_04047_));
 sky130_fd_sc_hd__and4_1 _10981_ (.A(_06416_),
    .B(_00438_),
    .C(net109),
    .D(_02164_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_2 _10982_ (.A(_04047_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__and2_2 _10983_ (.A(_03455_),
    .B(_03457_),
    .X(_04050_));
 sky130_fd_sc_hd__xnor2_4 _10984_ (.A(_04049_),
    .B(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__o21ba_2 _10985_ (.A1(_03453_),
    .A2(_03460_),
    .B1_N(_03459_),
    .X(_04053_));
 sky130_fd_sc_hd__xnor2_4 _10986_ (.A(_04052_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__xor2_4 _10987_ (.A(_04046_),
    .B(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__a21oi_2 _10988_ (.A1(_03476_),
    .A2(_03465_),
    .B1(_03464_),
    .Y(_04056_));
 sky130_fd_sc_hd__xnor2_4 _10989_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__xnor2_4 _10990_ (.A(_04037_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand3_1 _10991_ (.A(_03487_),
    .B(_03501_),
    .C(_03503_),
    .Y(_04059_));
 sky130_fd_sc_hd__a21o_1 _10992_ (.A1(_03530_),
    .A2(_03549_),
    .B1(_03548_),
    .X(_04060_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_03496_),
    .B(_03500_),
    .Y(_04061_));
 sky130_fd_sc_hd__and2_1 _10994_ (.A(_02906_),
    .B(_03528_),
    .X(_04063_));
 sky130_fd_sc_hd__a21o_1 _10995_ (.A1(_03525_),
    .A2(_03529_),
    .B1(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__a22o_1 _10996_ (.A1(net134),
    .A2(net178),
    .B1(net145),
    .B2(net177),
    .X(_04065_));
 sky130_fd_sc_hd__nand4_1 _10997_ (.A(_00453_),
    .B(net134),
    .C(net178),
    .D(net145),
    .Y(_04066_));
 sky130_fd_sc_hd__and2_1 _10998_ (.A(net123),
    .B(net180),
    .X(_04067_));
 sky130_fd_sc_hd__a21o_1 _10999_ (.A1(_04065_),
    .A2(_04066_),
    .B1(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__nand3_1 _11000_ (.A(_04065_),
    .B(_04066_),
    .C(_04067_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21bo_1 _11001_ (.A1(_03489_),
    .A2(_03492_),
    .B1_N(_03490_),
    .X(_04070_));
 sky130_fd_sc_hd__nand3_1 _11002_ (.A(_04068_),
    .B(_04069_),
    .C(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__a21o_1 _11003_ (.A1(_04068_),
    .A2(_04069_),
    .B1(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__a22o_1 _11004_ (.A1(_00059_),
    .A2(_03499_),
    .B1(_04071_),
    .B2(_04072_),
    .X(_04074_));
 sky130_fd_sc_hd__nand4_1 _11005_ (.A(_00059_),
    .B(_03499_),
    .C(_04071_),
    .D(_04072_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand3_1 _11006_ (.A(_04064_),
    .B(_04074_),
    .C(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__a21o_1 _11007_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04064_),
    .X(_04077_));
 sky130_fd_sc_hd__nand3_1 _11008_ (.A(_04061_),
    .B(_04076_),
    .C(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__a21o_1 _11009_ (.A1(_04076_),
    .A2(_04077_),
    .B1(_04061_),
    .X(_04079_));
 sky130_fd_sc_hd__and3_1 _11010_ (.A(_04060_),
    .B(_04078_),
    .C(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__a21oi_1 _11011_ (.A1(_04078_),
    .A2(_04079_),
    .B1(_04060_),
    .Y(_04081_));
 sky130_fd_sc_hd__a211o_2 _11012_ (.A1(_03501_),
    .A2(_04059_),
    .B1(_04080_),
    .C1(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__o211ai_2 _11013_ (.A1(_04080_),
    .A2(_04081_),
    .B1(_03501_),
    .C1(_04059_),
    .Y(_04083_));
 sky130_fd_sc_hd__o211a_1 _11014_ (.A1(_03506_),
    .A2(_03508_),
    .B1(_04082_),
    .C1(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__a211oi_2 _11015_ (.A1(_04082_),
    .A2(_04083_),
    .B1(_03506_),
    .C1(_03508_),
    .Y(_04086_));
 sky130_fd_sc_hd__or3_1 _11016_ (.A(_04058_),
    .B(_04085_),
    .C(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__o21ai_1 _11017_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_04058_),
    .Y(_04088_));
 sky130_fd_sc_hd__o211a_1 _11018_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04087_),
    .C1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a211o_1 _11019_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04024_),
    .C1(_04025_),
    .X(_04090_));
 sky130_fd_sc_hd__or2b_2 _11020_ (.A(_04089_),
    .B_N(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__xnor2_4 _11021_ (.A(_04023_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__nor2_1 _11022_ (.A(_03562_),
    .B(_03564_),
    .Y(_04093_));
 sky130_fd_sc_hd__a21o_2 _11023_ (.A1(_03551_),
    .A2(_03565_),
    .B1(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__nor2_1 _11024_ (.A(_03572_),
    .B(_03598_),
    .Y(_04096_));
 sky130_fd_sc_hd__a21o_2 _11025_ (.A1(_03571_),
    .A2(_03599_),
    .B1(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__a22o_1 _11026_ (.A1(_00489_),
    .A2(net197),
    .B1(net198),
    .B2(_00049_),
    .X(_04098_));
 sky130_fd_sc_hd__and4_2 _11027_ (.A(_00047_),
    .B(net186),
    .C(net197),
    .D(net198),
    .X(_04099_));
 sky130_fd_sc_hd__inv_2 _11028_ (.A(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__and2_1 _11029_ (.A(_04098_),
    .B(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__nand4_1 _11030_ (.A(_00058_),
    .B(_00481_),
    .C(net188),
    .D(net189),
    .Y(_04102_));
 sky130_fd_sc_hd__a22o_1 _11031_ (.A1(_00480_),
    .A2(net188),
    .B1(net189),
    .B2(_00989_),
    .X(_04103_));
 sky130_fd_sc_hd__and2_1 _11032_ (.A(_01002_),
    .B(net196),
    .X(_04104_));
 sky130_fd_sc_hd__a21o_1 _11033_ (.A1(_04102_),
    .A2(_04103_),
    .B1(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__nand3_1 _11034_ (.A(_04102_),
    .B(_04103_),
    .C(_04104_),
    .Y(_04107_));
 sky130_fd_sc_hd__a21bo_1 _11035_ (.A1(_03537_),
    .A2(_03539_),
    .B1_N(_03538_),
    .X(_04108_));
 sky130_fd_sc_hd__nand3_2 _11036_ (.A(_04105_),
    .B(_04107_),
    .C(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__a21o_1 _11037_ (.A1(_04105_),
    .A2(_04107_),
    .B1(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__nand3_2 _11038_ (.A(_04101_),
    .B(_04109_),
    .C(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21o_1 _11039_ (.A1(_04109_),
    .A2(_04110_),
    .B1(_04101_),
    .X(_04112_));
 sky130_fd_sc_hd__a21bo_1 _11040_ (.A1(_03533_),
    .A2(_03543_),
    .B1_N(_03542_),
    .X(_04113_));
 sky130_fd_sc_hd__and3_1 _11041_ (.A(_04111_),
    .B(_04112_),
    .C(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__a21o_1 _11042_ (.A1(_04111_),
    .A2(_04112_),
    .B1(_04113_),
    .X(_04115_));
 sky130_fd_sc_hd__and2b_1 _11043_ (.A_N(_04114_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _11044_ (.A(_05202_),
    .B(_01563_),
    .Y(_04118_));
 sky130_fd_sc_hd__and3_1 _11045_ (.A(_00062_),
    .B(_02215_),
    .C(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__xor2_4 _11046_ (.A(_03532_),
    .B(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__xnor2_4 _11047_ (.A(_04116_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a21o_1 _11048_ (.A1(_03577_),
    .A2(_03587_),
    .B1(_03586_),
    .X(_04122_));
 sky130_fd_sc_hd__buf_2 _11049_ (.A(net233),
    .X(_04123_));
 sky130_fd_sc_hd__and3_1 _11050_ (.A(_04752_),
    .B(_04123_),
    .C(_03575_),
    .X(_04124_));
 sky130_fd_sc_hd__nor2_1 _11051_ (.A(_03574_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__xnor2_2 _11052_ (.A(_04122_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__or2b_1 _11053_ (.A(_03556_),
    .B_N(_03558_),
    .X(_04127_));
 sky130_fd_sc_hd__and3_1 _11054_ (.A(_05093_),
    .B(_02239_),
    .C(_04127_),
    .X(_04129_));
 sky130_fd_sc_hd__xnor2_2 _11055_ (.A(_04126_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__and2_1 _11056_ (.A(_03555_),
    .B(_03560_),
    .X(_04131_));
 sky130_fd_sc_hd__a21oi_2 _11057_ (.A1(_03553_),
    .A2(_03561_),
    .B1(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__xor2_2 _11058_ (.A(_04130_),
    .B(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__xnor2_4 _11059_ (.A(_04121_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__xnor2_4 _11060_ (.A(_04097_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xnor2_4 _11061_ (.A(_04094_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__or2b_1 _11062_ (.A(_03594_),
    .B_N(_03596_),
    .X(_04137_));
 sky130_fd_sc_hd__o21ai_4 _11063_ (.A1(_03589_),
    .A2(_03597_),
    .B1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a21oi_1 _11064_ (.A1(_03602_),
    .A2(_03617_),
    .B1(_03616_),
    .Y(_04140_));
 sky130_fd_sc_hd__a22oi_1 _11065_ (.A1(net222),
    .A2(net231),
    .B1(_01603_),
    .B2(net221),
    .Y(_04141_));
 sky130_fd_sc_hd__and4_1 _11066_ (.A(net221),
    .B(net222),
    .C(net231),
    .D(net232),
    .X(_04142_));
 sky130_fd_sc_hd__or2_1 _11067_ (.A(_04141_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(_00080_),
    .B(_04123_),
    .Y(_04144_));
 sky130_fd_sc_hd__xnor2_2 _11069_ (.A(_04143_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a22oi_1 _11070_ (.A1(_00516_),
    .A2(_01617_),
    .B1(_03580_),
    .B2(_00086_),
    .Y(_04146_));
 sky130_fd_sc_hd__and4_1 _11071_ (.A(_00086_),
    .B(net230),
    .C(net224),
    .D(_03580_),
    .X(_04147_));
 sky130_fd_sc_hd__nor2_1 _11072_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__a21bo_1 _11073_ (.A1(_03578_),
    .A2(_03582_),
    .B1_N(_03581_),
    .X(_04149_));
 sky130_fd_sc_hd__xor2_2 _11074_ (.A(_04148_),
    .B(_04149_),
    .X(_04151_));
 sky130_fd_sc_hd__xnor2_2 _11075_ (.A(_04145_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__a31o_1 _11076_ (.A1(_00107_),
    .A2(_01629_),
    .A3(_03606_),
    .B1(_03605_),
    .X(_04153_));
 sky130_fd_sc_hd__buf_2 _11077_ (.A(net49),
    .X(_04154_));
 sky130_fd_sc_hd__nand2_1 _11078_ (.A(_00107_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__xor2_1 _11079_ (.A(_04153_),
    .B(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__and3_1 _11080_ (.A(_04906_),
    .B(_04154_),
    .C(_03591_),
    .X(_04157_));
 sky130_fd_sc_hd__a21oi_1 _11081_ (.A1(_02969_),
    .A2(_03593_),
    .B1(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__xor2_1 _11082_ (.A(_04156_),
    .B(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__xnor2_1 _11083_ (.A(_04152_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__nor2_1 _11084_ (.A(_04140_),
    .B(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__and2_1 _11085_ (.A(_04140_),
    .B(_04160_),
    .X(_04163_));
 sky130_fd_sc_hd__nor2_2 _11086_ (.A(_04162_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__xor2_4 _11087_ (.A(_04138_),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__and2b_1 _11088_ (.A_N(_03608_),
    .B(_03614_),
    .X(_04166_));
 sky130_fd_sc_hd__a21o_2 _11089_ (.A1(_03611_),
    .A2(_03613_),
    .B1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__and2_1 _11090_ (.A(_03621_),
    .B(_03625_),
    .X(_04168_));
 sky130_fd_sc_hd__a22oi_1 _11091_ (.A1(_01068_),
    .A2(_01051_),
    .B1(_01653_),
    .B2(_00530_),
    .Y(_04169_));
 sky130_fd_sc_hd__and4_1 _11092_ (.A(net46),
    .B(net38),
    .C(net47),
    .D(net39),
    .X(_04170_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(_00543_),
    .B(net48),
    .Y(_04173_));
 sky130_fd_sc_hd__xor2_1 _11095_ (.A(_04171_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__nand2_1 _11096_ (.A(_04862_),
    .B(_01653_),
    .Y(_04175_));
 sky130_fd_sc_hd__and3_1 _11097_ (.A(_00097_),
    .B(_02329_),
    .C(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__xnor2_1 _11098_ (.A(_04174_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__o21a_1 _11099_ (.A1(_04168_),
    .A2(_03628_),
    .B1(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__or3_1 _11100_ (.A(_04168_),
    .B(_03628_),
    .C(_04177_),
    .X(_04179_));
 sky130_fd_sc_hd__or2b_2 _11101_ (.A(_04178_),
    .B_N(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__xnor2_4 _11102_ (.A(_04167_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__a22o_1 _11103_ (.A1(_00544_),
    .A2(_01667_),
    .B1(net234),
    .B2(_00109_),
    .X(_04182_));
 sky130_fd_sc_hd__nand4_1 _11104_ (.A(_00109_),
    .B(_00544_),
    .C(_01667_),
    .D(_03019_),
    .Y(_04184_));
 sky130_fd_sc_hd__and2_1 _11105_ (.A(_01666_),
    .B(net45),
    .X(_04185_));
 sky130_fd_sc_hd__a21o_1 _11106_ (.A1(_04182_),
    .A2(_04184_),
    .B1(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__nand3_1 _11107_ (.A(_04182_),
    .B(_04184_),
    .C(_04185_),
    .Y(_04187_));
 sky130_fd_sc_hd__o211a_1 _11108_ (.A1(_03022_),
    .A2(_03639_),
    .B1(_04186_),
    .C1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__a211o_1 _11109_ (.A1(_04186_),
    .A2(_04187_),
    .B1(_03022_),
    .C1(_03639_),
    .X(_04189_));
 sky130_fd_sc_hd__or2b_2 _11110_ (.A(_04188_),
    .B_N(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__a21bo_2 _11111_ (.A1(_03630_),
    .A2(_03632_),
    .B1_N(_03631_),
    .X(_04191_));
 sky130_fd_sc_hd__a22oi_1 _11112_ (.A1(_00550_),
    .A2(_01652_),
    .B1(_03006_),
    .B2(_00549_),
    .Y(_04192_));
 sky130_fd_sc_hd__and4_2 _11113_ (.A(_00549_),
    .B(_00550_),
    .C(net56),
    .D(_03006_),
    .X(_04193_));
 sky130_fd_sc_hd__nor2_2 _11114_ (.A(_04192_),
    .B(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__xor2_4 _11115_ (.A(_04191_),
    .B(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__xor2_4 _11116_ (.A(_03624_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__xnor2_4 _11117_ (.A(_04190_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__and2b_1 _11118_ (.A_N(_03642_),
    .B(_03640_),
    .X(_04199_));
 sky130_fd_sc_hd__a21o_1 _11119_ (.A1(_03629_),
    .A2(_03643_),
    .B1(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__xor2_4 _11120_ (.A(_04198_),
    .B(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__xnor2_4 _11121_ (.A(_04181_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(_03644_),
    .B(_03647_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21bo_1 _11123_ (.A1(_03619_),
    .A2(_03648_),
    .B1_N(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__xnor2_4 _11124_ (.A(_04202_),
    .B(_04204_),
    .Y(_04206_));
 sky130_fd_sc_hd__xnor2_4 _11125_ (.A(_04165_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__or2b_1 _11126_ (.A(_03651_),
    .B_N(_03649_),
    .X(_04208_));
 sky130_fd_sc_hd__a21bo_2 _11127_ (.A1(_03600_),
    .A2(_03652_),
    .B1_N(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__xnor2_4 _11128_ (.A(_04207_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_4 _11129_ (.A(_04136_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__and2b_1 _11130_ (.A_N(_03653_),
    .B(_03655_),
    .X(_04212_));
 sky130_fd_sc_hd__a21oi_4 _11131_ (.A1(_03569_),
    .A2(_03657_),
    .B1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__xor2_4 _11132_ (.A(_04211_),
    .B(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__xnor2_4 _11133_ (.A(_04092_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nor2_1 _11134_ (.A(_03658_),
    .B(_03660_),
    .Y(_04217_));
 sky130_fd_sc_hd__a21oi_2 _11135_ (.A1(_03519_),
    .A2(_03661_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__xor2_4 _11136_ (.A(_04215_),
    .B(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__xnor2_4 _11137_ (.A(_04022_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _11138_ (.A(_03662_),
    .B(_03664_),
    .Y(_04221_));
 sky130_fd_sc_hd__a21oi_4 _11139_ (.A1(_03431_),
    .A2(_03665_),
    .B1(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__xor2_4 _11140_ (.A(_04220_),
    .B(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__xnor2_4 _11141_ (.A(_03915_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__nor2_1 _11142_ (.A(_03666_),
    .B(_03669_),
    .Y(_04225_));
 sky130_fd_sc_hd__a21oi_4 _11143_ (.A1(_03316_),
    .A2(_03670_),
    .B1(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__xor2_2 _11144_ (.A(_04224_),
    .B(_04226_),
    .X(_04228_));
 sky130_fd_sc_hd__xnor2_2 _11145_ (.A(_03739_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nor2_1 _11146_ (.A(_03671_),
    .B(_03673_),
    .Y(_04230_));
 sky130_fd_sc_hd__a21oi_2 _11147_ (.A1(_03125_),
    .A2(_03674_),
    .B1(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__xor2_2 _11148_ (.A(_04229_),
    .B(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__xnor2_2 _11149_ (.A(_03695_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__nor2_1 _11150_ (.A(_03675_),
    .B(_03677_),
    .Y(_04234_));
 sky130_fd_sc_hd__a21oi_2 _11151_ (.A1(_03079_),
    .A2(_03679_),
    .B1(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__xor2_2 _11152_ (.A(_04233_),
    .B(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__and2_1 _11153_ (.A(_03061_),
    .B(_03683_),
    .X(_04237_));
 sky130_fd_sc_hd__a21o_1 _11154_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03680_),
    .X(_04239_));
 sky130_fd_sc_hd__a21oi_1 _11155_ (.A1(_03074_),
    .A2(_04239_),
    .B1(_03682_),
    .Y(_04240_));
 sky130_fd_sc_hd__a21o_1 _11156_ (.A1(_03065_),
    .A2(_04237_),
    .B1(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__xor2_1 _11157_ (.A(_04236_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_1 _11158_ (.A(net259),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__or2_1 _11159_ (.A(net259),
    .B(_04242_),
    .X(_04244_));
 sky130_fd_sc_hd__and2_1 _11160_ (.A(_04243_),
    .B(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__a21o_1 _11161_ (.A1(_03691_),
    .A2(_03692_),
    .B1(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__nand3_1 _11162_ (.A(_03691_),
    .B(_03692_),
    .C(_04245_),
    .Y(_04247_));
 sky130_fd_sc_hd__and3_1 _11163_ (.A(_02185_),
    .B(_04246_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_04248_),
    .X(_00010_));
 sky130_fd_sc_hd__nor2_1 _11165_ (.A(_04233_),
    .B(_04235_),
    .Y(_04250_));
 sky130_fd_sc_hd__a21oi_1 _11166_ (.A1(_04236_),
    .A2(_04241_),
    .B1(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__nor2_1 _11167_ (.A(_04229_),
    .B(_04231_),
    .Y(_04252_));
 sky130_fd_sc_hd__a21oi_2 _11168_ (.A1(_03695_),
    .A2(_04232_),
    .B1(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__or2b_1 _11169_ (.A(_03737_),
    .B_N(_03700_),
    .X(_04254_));
 sky130_fd_sc_hd__or2b_1 _11170_ (.A(_03738_),
    .B_N(_03697_),
    .X(_04255_));
 sky130_fd_sc_hd__nand2_1 _11171_ (.A(_04254_),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__or2b_1 _11172_ (.A(_03703_),
    .B_N(_03735_),
    .X(_04257_));
 sky130_fd_sc_hd__a21bo_2 _11173_ (.A1(_03702_),
    .A2(_03736_),
    .B1_N(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__and2b_1 _11174_ (.A_N(_03913_),
    .B(_03741_),
    .X(_04260_));
 sky130_fd_sc_hd__a21o_2 _11175_ (.A1(_03740_),
    .A2(_03914_),
    .B1(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__and2b_1 _11176_ (.A_N(_03704_),
    .B(_03734_),
    .X(_04262_));
 sky130_fd_sc_hd__nor2_2 _11177_ (.A(_03731_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__a21o_2 _11178_ (.A1(_03768_),
    .A2(_03847_),
    .B1(_03845_),
    .X(_04264_));
 sky130_fd_sc_hd__a31o_2 _11179_ (.A1(_06243_),
    .A2(_01754_),
    .A3(_03728_),
    .B1(_03726_),
    .X(_04265_));
 sky130_fd_sc_hd__or2b_1 _11180_ (.A(_03746_),
    .B_N(_03766_),
    .X(_04266_));
 sky130_fd_sc_hd__or2b_1 _11181_ (.A(_03744_),
    .B_N(_03767_),
    .X(_04267_));
 sky130_fd_sc_hd__o21a_1 _11182_ (.A1(_03723_),
    .A2(_03724_),
    .B1(_03720_),
    .X(_04268_));
 sky130_fd_sc_hd__a22o_1 _11183_ (.A1(_00617_),
    .A2(_01188_),
    .B1(_02464_),
    .B2(_00171_),
    .X(_04269_));
 sky130_fd_sc_hd__nand3_1 _11184_ (.A(_00617_),
    .B(_02464_),
    .C(_03709_),
    .Y(_04271_));
 sky130_fd_sc_hd__or2_1 _11185_ (.A(_03712_),
    .B(_03714_),
    .X(_04272_));
 sky130_fd_sc_hd__and3_1 _11186_ (.A(_04269_),
    .B(_04271_),
    .C(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a21oi_1 _11187_ (.A1(_04269_),
    .A2(_04271_),
    .B1(_04272_),
    .Y(_04274_));
 sky130_fd_sc_hd__nor2_1 _11188_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_1 _11189_ (.A(_03717_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(_01777_),
    .B(_01157_),
    .Y(_04277_));
 sky130_fd_sc_hd__xnor2_1 _11191_ (.A(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__and2b_1 _11192_ (.A_N(_04268_),
    .B(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__and2b_1 _11193_ (.A_N(_04278_),
    .B(_04268_),
    .X(_04280_));
 sky130_fd_sc_hd__nor2_1 _11194_ (.A(_04279_),
    .B(_04280_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_1 _11195_ (.A(_00270_),
    .B(_01754_),
    .Y(_04283_));
 sky130_fd_sc_hd__xor2_1 _11196_ (.A(_04282_),
    .B(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__a21oi_1 _11197_ (.A1(_04266_),
    .A2(_04267_),
    .B1(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__and3_1 _11198_ (.A(_04266_),
    .B(_04267_),
    .C(_04284_),
    .X(_04286_));
 sky130_fd_sc_hd__nor2_2 _11199_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__xnor2_4 _11200_ (.A(_04265_),
    .B(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__xnor2_2 _11201_ (.A(_04264_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__xnor2_2 _11202_ (.A(_04263_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_2 _11203_ (.A(_04261_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__xnor2_2 _11204_ (.A(_04258_),
    .B(_04291_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21o_2 _11205_ (.A1(_03848_),
    .A2(_03912_),
    .B1(_03910_),
    .X(_04294_));
 sky130_fd_sc_hd__a21o_2 _11206_ (.A1(_03917_),
    .A2(_04020_),
    .B1(_04019_),
    .X(_04295_));
 sky130_fd_sc_hd__or2b_1 _11207_ (.A(_03748_),
    .B_N(_03763_),
    .X(_04296_));
 sky130_fd_sc_hd__or2b_1 _11208_ (.A(_03747_),
    .B_N(_03764_),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _11209_ (.A(_04296_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__a21o_1 _11210_ (.A1(_03794_),
    .A2(_03810_),
    .B1(_03807_),
    .X(_04299_));
 sky130_fd_sc_hd__and2b_1 _11211_ (.A_N(_03750_),
    .B(_03762_),
    .X(_04300_));
 sky130_fd_sc_hd__a31oi_2 _11212_ (.A1(_03751_),
    .A2(_03759_),
    .A3(_03760_),
    .B1(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _11213_ (.A1(_03777_),
    .A2(_03792_),
    .B1(_03791_),
    .Y(_04302_));
 sky130_fd_sc_hd__a22o_1 _11214_ (.A1(net29),
    .A2(_01217_),
    .B1(_01181_),
    .B2(net20),
    .X(_04304_));
 sky130_fd_sc_hd__inv_2 _11215_ (.A(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__and4_1 _11216_ (.A(_00706_),
    .B(_00647_),
    .C(_01217_),
    .D(_01181_),
    .X(_04306_));
 sky130_fd_sc_hd__o2bb2a_1 _11217_ (.A1_N(_00239_),
    .A2_N(_01784_),
    .B1(_04305_),
    .B2(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__and4b_1 _11218_ (.A_N(_04306_),
    .B(_01784_),
    .C(_00239_),
    .D(_04304_),
    .X(_04308_));
 sky130_fd_sc_hd__a41o_1 _11219_ (.A1(_00239_),
    .A2(_00706_),
    .A3(_00647_),
    .A4(_01181_),
    .B1(_03756_),
    .X(_04309_));
 sky130_fd_sc_hd__or3b_2 _11220_ (.A(_04307_),
    .B(_04308_),
    .C_N(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__o21bai_1 _11221_ (.A1(_04307_),
    .A2(_04308_),
    .B1_N(_04309_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _11222_ (.A(_04310_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__xor2_1 _11223_ (.A(_03774_),
    .B(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__xnor2_1 _11224_ (.A(_03759_),
    .B(_04313_),
    .Y(_04315_));
 sky130_fd_sc_hd__xnor2_1 _11225_ (.A(_04302_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__xnor2_1 _11226_ (.A(_04301_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__xor2_1 _11227_ (.A(_04299_),
    .B(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__xnor2_1 _11228_ (.A(_04298_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a22o_1 _11229_ (.A1(_00703_),
    .A2(net92),
    .B1(_01858_),
    .B2(_00238_),
    .X(_04320_));
 sky130_fd_sc_hd__and4_1 _11230_ (.A(net98),
    .B(net99),
    .C(net92),
    .D(net93),
    .X(_04321_));
 sky130_fd_sc_hd__inv_2 _11231_ (.A(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__and4_1 _11232_ (.A(_00672_),
    .B(_01835_),
    .C(_04320_),
    .D(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__a22oi_1 _11233_ (.A1(_00672_),
    .A2(_01835_),
    .B1(_04320_),
    .B2(_04322_),
    .Y(_04324_));
 sky130_fd_sc_hd__nor2_1 _11234_ (.A(_04323_),
    .B(_04324_),
    .Y(_04326_));
 sky130_fd_sc_hd__o21ba_1 _11235_ (.A1(_03780_),
    .A2(_03783_),
    .B1_N(_03781_),
    .X(_04327_));
 sky130_fd_sc_hd__xnor2_2 _11236_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(_00200_),
    .B(_03180_),
    .Y(_04329_));
 sky130_fd_sc_hd__xor2_2 _11238_ (.A(_04328_),
    .B(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__a31o_1 _11239_ (.A1(_06284_),
    .A2(_03180_),
    .A3(_03788_),
    .B1(_03785_),
    .X(_04331_));
 sky130_fd_sc_hd__xnor2_2 _11240_ (.A(_04330_),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _11241_ (.A(_06264_),
    .B(_01217_),
    .Y(_04333_));
 sky130_fd_sc_hd__and3_1 _11242_ (.A(_00250_),
    .B(_02498_),
    .C(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__xnor2_2 _11243_ (.A(_04332_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21a_1 _11244_ (.A1(_03797_),
    .A2(_03801_),
    .B1(_03803_),
    .X(_04337_));
 sky130_fd_sc_hd__a21oi_1 _11245_ (.A1(_06134_),
    .A2(_01251_),
    .B1(_03212_),
    .Y(_04338_));
 sky130_fd_sc_hd__nor2_1 _11246_ (.A(_03799_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__xnor2_1 _11247_ (.A(_03817_),
    .B(_03826_),
    .Y(_04340_));
 sky130_fd_sc_hd__o31ai_2 _11248_ (.A1(_03816_),
    .A2(_03817_),
    .A3(_03828_),
    .B1(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__xor2_1 _11249_ (.A(_04339_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__or2b_1 _11250_ (.A(_04337_),
    .B_N(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__or2b_1 _11251_ (.A(_04342_),
    .B_N(_04337_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_1 _11252_ (.A(_04343_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__xor2_2 _11253_ (.A(_04335_),
    .B(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _11254_ (.A(_03830_),
    .B(_03833_),
    .Y(_04348_));
 sky130_fd_sc_hd__o21ai_4 _11255_ (.A1(_03829_),
    .A2(_03834_),
    .B1(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__a21bo_2 _11256_ (.A1(_03858_),
    .A2(_03874_),
    .B1_N(_03873_),
    .X(_04350_));
 sky130_fd_sc_hd__a32o_1 _11257_ (.A1(_06311_),
    .A2(_02592_),
    .A3(_03862_),
    .B1(_03861_),
    .B2(_00749_),
    .X(_04351_));
 sky130_fd_sc_hd__a22o_1 _11258_ (.A1(_00677_),
    .A2(net137),
    .B1(net138),
    .B2(_00210_),
    .X(_04352_));
 sky130_fd_sc_hd__and4_1 _11259_ (.A(_00210_),
    .B(_00677_),
    .C(net137),
    .D(net138),
    .X(_04353_));
 sky130_fd_sc_hd__inv_2 _11260_ (.A(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__and2_1 _11261_ (.A(_04352_),
    .B(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__a22oi_1 _11262_ (.A1(net136),
    .A2(net128),
    .B1(net129),
    .B2(_00201_),
    .Y(_04356_));
 sky130_fd_sc_hd__and4_1 _11263_ (.A(net135),
    .B(net136),
    .C(net128),
    .D(net129),
    .X(_04357_));
 sky130_fd_sc_hd__nor2_1 _11264_ (.A(_04356_),
    .B(_04357_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21bo_1 _11265_ (.A1(_03819_),
    .A2(_03822_),
    .B1_N(_03821_),
    .X(_04360_));
 sky130_fd_sc_hd__nand2_1 _11266_ (.A(_04359_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__or2_1 _11267_ (.A(_04359_),
    .B(_04360_),
    .X(_04362_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(_04361_),
    .B(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__xor2_1 _11269_ (.A(_04355_),
    .B(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__and2_2 _11270_ (.A(_04351_),
    .B(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _11271_ (.A(_04351_),
    .B(_04364_),
    .Y(_04366_));
 sky130_fd_sc_hd__or2_2 _11272_ (.A(_04365_),
    .B(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__xnor2_4 _11273_ (.A(_04350_),
    .B(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__xnor2_4 _11274_ (.A(_04349_),
    .B(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__and2_1 _11275_ (.A(_03815_),
    .B(_03835_),
    .X(_04371_));
 sky130_fd_sc_hd__a21o_2 _11276_ (.A1(_03814_),
    .A2(_03836_),
    .B1(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__xnor2_4 _11277_ (.A(_04370_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__xnor2_2 _11278_ (.A(_04346_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__o21a_1 _11279_ (.A1(_03811_),
    .A2(_03843_),
    .B1(_03840_),
    .X(_04375_));
 sky130_fd_sc_hd__xnor2_1 _11280_ (.A(_04374_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__or2_2 _11281_ (.A(_04319_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__nand2_1 _11282_ (.A(_04319_),
    .B(_04376_),
    .Y(_04378_));
 sky130_fd_sc_hd__and2_2 _11283_ (.A(_04377_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__or2b_1 _11284_ (.A(_03903_),
    .B_N(_03855_),
    .X(_04381_));
 sky130_fd_sc_hd__a21bo_1 _11285_ (.A1(_03857_),
    .A2(_03902_),
    .B1_N(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__or2b_1 _11286_ (.A(_03978_),
    .B_N(_03976_),
    .X(_04383_));
 sky130_fd_sc_hd__a21boi_2 _11287_ (.A1(_03936_),
    .A2(_03979_),
    .B1_N(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__and2b_1 _11288_ (.A_N(_03900_),
    .B(_03896_),
    .X(_04385_));
 sky130_fd_sc_hd__a21o_1 _11289_ (.A1(_03878_),
    .A2(_03901_),
    .B1(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__and2_1 _11290_ (.A(_03922_),
    .B(_03934_),
    .X(_04387_));
 sky130_fd_sc_hd__a21o_2 _11291_ (.A1(_03921_),
    .A2(_03935_),
    .B1(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__and3_1 _11292_ (.A(_00774_),
    .B(net153),
    .C(_01288_),
    .X(_04389_));
 sky130_fd_sc_hd__a22o_1 _11293_ (.A1(net153),
    .A2(net146),
    .B1(_01288_),
    .B2(_00774_),
    .X(_04390_));
 sky130_fd_sc_hd__a21bo_1 _11294_ (.A1(_01309_),
    .A2(_04389_),
    .B1_N(_04390_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _11295_ (.A(_00291_),
    .B(_02592_),
    .Y(_04393_));
 sky130_fd_sc_hd__xnor2_1 _11296_ (.A(_04392_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _11297_ (.A(_06319_),
    .B(_01309_),
    .Y(_04395_));
 sky130_fd_sc_hd__and3_1 _11298_ (.A(_01293_),
    .B(_02615_),
    .C(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__xnor2_1 _11299_ (.A(_04394_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__xnor2_1 _11300_ (.A(_03881_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a32o_1 _11301_ (.A1(_03867_),
    .A2(_03868_),
    .A3(_03870_),
    .B1(_03871_),
    .B2(_03866_),
    .X(_04399_));
 sky130_fd_sc_hd__and2b_1 _11302_ (.A_N(_04398_),
    .B(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__and2b_1 _11303_ (.A_N(_04399_),
    .B(_04398_),
    .X(_04401_));
 sky130_fd_sc_hd__nor2_1 _11304_ (.A(_04400_),
    .B(_04401_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _11305_ (.A(_03885_),
    .B(_03888_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _11306_ (.A(_00343_),
    .B(net216),
    .Y(_04405_));
 sky130_fd_sc_hd__xor2_1 _11307_ (.A(_04404_),
    .B(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__a22oi_1 _11308_ (.A1(_00757_),
    .A2(_01365_),
    .B1(_01986_),
    .B2(_00297_),
    .Y(_04407_));
 sky130_fd_sc_hd__and4_1 _11309_ (.A(_00297_),
    .B(net214),
    .C(net206),
    .D(net207),
    .X(_04408_));
 sky130_fd_sc_hd__nor2_1 _11310_ (.A(_04407_),
    .B(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(_00810_),
    .B(_02626_),
    .Y(_04410_));
 sky130_fd_sc_hd__xnor2_1 _11312_ (.A(_04409_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__a31o_1 _11313_ (.A1(_03887_),
    .A2(_03888_),
    .A3(_03891_),
    .B1(_03292_),
    .X(_04412_));
 sky130_fd_sc_hd__xnor2_1 _11314_ (.A(_04411_),
    .B(_04412_),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_1 _11315_ (.A(_04406_),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__and2_1 _11316_ (.A(_04406_),
    .B(_04414_),
    .X(_04416_));
 sky130_fd_sc_hd__or2_1 _11317_ (.A(_04415_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_1 _11318_ (.A(_03892_),
    .B(_03894_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21o_1 _11319_ (.A1(_03883_),
    .A2(_03895_),
    .B1(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__xnor2_2 _11320_ (.A(_04417_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__xor2_2 _11321_ (.A(_04403_),
    .B(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__xnor2_2 _11322_ (.A(_04388_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__xor2_2 _11323_ (.A(_04386_),
    .B(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__xor2_2 _11324_ (.A(_04384_),
    .B(_04423_),
    .X(_04425_));
 sky130_fd_sc_hd__xnor2_1 _11325_ (.A(_04382_),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2_1 _11326_ (.A(_03852_),
    .B(_03904_),
    .Y(_04427_));
 sky130_fd_sc_hd__a21boi_2 _11327_ (.A1(_03850_),
    .A2(_03905_),
    .B1_N(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__nor2_1 _11328_ (.A(_04426_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_04426_),
    .B(_04428_),
    .Y(_04430_));
 sky130_fd_sc_hd__and2b_1 _11330_ (.A_N(_04429_),
    .B(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__xnor2_4 _11331_ (.A(_04379_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__xnor2_4 _11332_ (.A(_04295_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__xor2_4 _11333_ (.A(_04294_),
    .B(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(_04013_),
    .B(_04015_),
    .Y(_04436_));
 sky130_fd_sc_hd__a21o_2 _11335_ (.A1(_03980_),
    .A2(_04016_),
    .B1(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__a21oi_2 _11336_ (.A1(_04023_),
    .A2(_04090_),
    .B1(_04089_),
    .Y(_04438_));
 sky130_fd_sc_hd__and2b_1 _11337_ (.A_N(_03933_),
    .B(_03924_),
    .X(_04439_));
 sky130_fd_sc_hd__a21o_1 _11338_ (.A1(_03925_),
    .A2(_03932_),
    .B1(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__o21ba_1 _11339_ (.A1(_03943_),
    .A2(_03958_),
    .B1_N(_03957_),
    .X(_04441_));
 sky130_fd_sc_hd__a22oi_1 _11340_ (.A1(_01385_),
    .A2(_01367_),
    .B1(_01987_),
    .B2(_00834_),
    .Y(_04442_));
 sky130_fd_sc_hd__and4_1 _11341_ (.A(_00834_),
    .B(_01385_),
    .C(_01367_),
    .D(_01987_),
    .X(_04443_));
 sky130_fd_sc_hd__nor2_1 _11342_ (.A(_04442_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__o21ai_2 _11343_ (.A1(_03938_),
    .A2(_03942_),
    .B1(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__or3_1 _11344_ (.A(_03938_),
    .B(_03942_),
    .C(_04444_),
    .X(_04447_));
 sky130_fd_sc_hd__a21o_1 _11345_ (.A1(_04445_),
    .A2(_04447_),
    .B1(_03928_),
    .X(_04448_));
 sky130_fd_sc_hd__nand3_1 _11346_ (.A(_03928_),
    .B(_04445_),
    .C(_04447_),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_04448_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_03926_),
    .B(_03929_),
    .Y(_04451_));
 sky130_fd_sc_hd__o21ai_2 _11349_ (.A1(_03328_),
    .A2(_03931_),
    .B1(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__xor2_2 _11350_ (.A(_04450_),
    .B(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__xor2_2 _11351_ (.A(_04441_),
    .B(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__xor2_2 _11352_ (.A(_04440_),
    .B(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__a22oi_1 _11353_ (.A1(_00830_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_00366_),
    .Y(_04456_));
 sky130_fd_sc_hd__and4_1 _11354_ (.A(_00366_),
    .B(_00830_),
    .C(_02694_),
    .D(_02695_),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_1 _11355_ (.A(_04456_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__a22o_1 _11356_ (.A1(_00821_),
    .A2(_01410_),
    .B1(_01397_),
    .B2(_00850_),
    .X(_04460_));
 sky130_fd_sc_hd__nand4_1 _11357_ (.A(_00850_),
    .B(_00821_),
    .C(_01410_),
    .D(_01397_),
    .Y(_04461_));
 sky130_fd_sc_hd__a22o_1 _11358_ (.A1(_00357_),
    .A2(_02019_),
    .B1(_04460_),
    .B2(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__nand4_1 _11359_ (.A(_00357_),
    .B(_02019_),
    .C(_04460_),
    .D(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand3b_1 _11360_ (.A_N(_03965_),
    .B(_04462_),
    .C(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__a21bo_1 _11361_ (.A1(_04462_),
    .A2(_04463_),
    .B1_N(_03965_),
    .X(_04465_));
 sky130_fd_sc_hd__nand2_1 _11362_ (.A(_03948_),
    .B(_03950_),
    .Y(_04466_));
 sky130_fd_sc_hd__a21o_1 _11363_ (.A1(_04464_),
    .A2(_04465_),
    .B1(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__nand3_1 _11364_ (.A(_04464_),
    .B(_04465_),
    .C(_04466_),
    .Y(_04469_));
 sky130_fd_sc_hd__o21bai_2 _11365_ (.A1(_03945_),
    .A2(_03953_),
    .B1_N(_03951_),
    .Y(_04470_));
 sky130_fd_sc_hd__and3_1 _11366_ (.A(_04467_),
    .B(_04469_),
    .C(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__a21o_1 _11367_ (.A1(_04467_),
    .A2(_04469_),
    .B1(_04470_),
    .X(_04472_));
 sky130_fd_sc_hd__and2b_1 _11368_ (.A_N(_04471_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__xnor2_2 _11369_ (.A(_04459_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__a21oi_2 _11370_ (.A1(_03988_),
    .A2(_03994_),
    .B1(_03993_),
    .Y(_04475_));
 sky130_fd_sc_hd__and4_1 _11371_ (.A(_00387_),
    .B(_00822_),
    .C(_03967_),
    .D(_02731_),
    .X(_04476_));
 sky130_fd_sc_hd__a22oi_2 _11372_ (.A1(_00387_),
    .A2(_03967_),
    .B1(_02731_),
    .B2(_00822_),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_1 _11373_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__xnor2_2 _11374_ (.A(_04475_),
    .B(_04478_),
    .Y(_04480_));
 sky130_fd_sc_hd__xor2_2 _11375_ (.A(_03966_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__nand2_1 _11376_ (.A(_03962_),
    .B(_03969_),
    .Y(_04482_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(_03962_),
    .B(_03969_),
    .Y(_04483_));
 sky130_fd_sc_hd__a21o_1 _11378_ (.A1(_03961_),
    .A2(_04482_),
    .B1(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__xnor2_2 _11379_ (.A(_04481_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__xnor2_2 _11380_ (.A(_04474_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__or2b_1 _11381_ (.A(_03973_),
    .B_N(_03971_),
    .X(_04487_));
 sky130_fd_sc_hd__a21bo_1 _11382_ (.A1(_03960_),
    .A2(_03975_),
    .B1_N(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__xnor2_2 _11383_ (.A(_04486_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__xor2_1 _11384_ (.A(_04455_),
    .B(_04489_),
    .X(_04491_));
 sky130_fd_sc_hd__and2b_1 _11385_ (.A_N(_03987_),
    .B(_04009_),
    .X(_04492_));
 sky130_fd_sc_hd__a21o_1 _11386_ (.A1(_03986_),
    .A2(_04010_),
    .B1(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__and2b_1 _11387_ (.A_N(_04056_),
    .B(_04055_),
    .X(_04494_));
 sky130_fd_sc_hd__a21o_1 _11388_ (.A1(_04037_),
    .A2(_04057_),
    .B1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__and2_1 _11389_ (.A(_04004_),
    .B(_04006_),
    .X(_04496_));
 sky130_fd_sc_hd__a21o_1 _11390_ (.A1(_03997_),
    .A2(_04008_),
    .B1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nor2_1 _11391_ (.A(_04027_),
    .B(_04035_),
    .Y(_04498_));
 sky130_fd_sc_hd__a21o_1 _11392_ (.A1(_04026_),
    .A2(_04036_),
    .B1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__and3_1 _11393_ (.A(_00397_),
    .B(_00872_),
    .C(_01444_),
    .X(_04500_));
 sky130_fd_sc_hd__a22o_1 _11394_ (.A1(_00872_),
    .A2(net57),
    .B1(net58),
    .B2(_00397_),
    .X(_04502_));
 sky130_fd_sc_hd__a21bo_1 _11395_ (.A1(_02765_),
    .A2(_04500_),
    .B1_N(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__nand2_1 _11396_ (.A(_00879_),
    .B(_01434_),
    .Y(_04504_));
 sky130_fd_sc_hd__xor2_2 _11397_ (.A(_04503_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nand2_1 _11398_ (.A(_03990_),
    .B(_03992_),
    .Y(_04506_));
 sky130_fd_sc_hd__xnor2_2 _11399_ (.A(_04505_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21bai_2 _11400_ (.A1(_03998_),
    .A2(_04003_),
    .B1_N(_04002_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_1 _11401_ (.A(net72),
    .B(net84),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _11402_ (.A(net73),
    .B(_01443_),
    .Y(_04510_));
 sky130_fd_sc_hd__or2_1 _11403_ (.A(_04509_),
    .B(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__or2_1 _11404_ (.A(_03999_),
    .B(_04511_),
    .X(_04513_));
 sky130_fd_sc_hd__nand2_1 _11405_ (.A(_04509_),
    .B(_04510_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_03999_),
    .B(_04511_),
    .Y(_04515_));
 sky130_fd_sc_hd__and3_1 _11407_ (.A(_04513_),
    .B(_04514_),
    .C(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__xnor2_2 _11408_ (.A(_04508_),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__xor2_2 _11409_ (.A(_04507_),
    .B(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__xor2_2 _11410_ (.A(_04499_),
    .B(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_2 _11411_ (.A(_04497_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__xnor2_2 _11412_ (.A(_04495_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__xnor2_2 _11413_ (.A(_04493_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__and2b_1 _11414_ (.A_N(_04011_),
    .B(_03983_),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_2 _11415_ (.A1(_03982_),
    .A2(_04012_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__xor2_1 _11416_ (.A(_04522_),
    .B(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__xnor2_1 _11417_ (.A(_04491_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nor2_1 _11418_ (.A(_04438_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__nand2_1 _11419_ (.A(_04438_),
    .B(_04527_),
    .Y(_04529_));
 sky130_fd_sc_hd__and2b_1 _11420_ (.A_N(_04528_),
    .B(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__xor2_4 _11421_ (.A(_04437_),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__or2b_2 _11422_ (.A(_04085_),
    .B_N(_04087_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _11423_ (.A(_04097_),
    .B(_04134_),
    .Y(_04533_));
 sky130_fd_sc_hd__or2b_1 _11424_ (.A(_04135_),
    .B_N(_04094_),
    .X(_04535_));
 sky130_fd_sc_hd__and2b_1 _11425_ (.A_N(_04034_),
    .B(_04033_),
    .X(_04536_));
 sky130_fd_sc_hd__or3_1 _11426_ (.A(_04042_),
    .B(_04043_),
    .C(_04045_),
    .X(_04537_));
 sky130_fd_sc_hd__a22oi_2 _11427_ (.A1(_00937_),
    .A2(_01488_),
    .B1(_02799_),
    .B2(_00421_),
    .Y(_04538_));
 sky130_fd_sc_hd__and4_2 _11428_ (.A(_00421_),
    .B(net82),
    .C(_01488_),
    .D(net75),
    .X(_04539_));
 sky130_fd_sc_hd__or2_1 _11429_ (.A(_04538_),
    .B(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__a32o_1 _11430_ (.A1(_01487_),
    .A2(_00937_),
    .A3(_04030_),
    .B1(_04028_),
    .B2(_02799_),
    .X(_04541_));
 sky130_fd_sc_hd__xnor2_1 _11431_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__xnor2_1 _11432_ (.A(_04537_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _11433_ (.A(_04536_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(_04536_),
    .B(_04543_),
    .X(_04546_));
 sky130_fd_sc_hd__nor2_2 _11435_ (.A(_04544_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__a22o_1 _11436_ (.A1(_00910_),
    .A2(_01520_),
    .B1(_01484_),
    .B2(_00956_),
    .X(_04548_));
 sky130_fd_sc_hd__nand4_2 _11437_ (.A(_00956_),
    .B(_00910_),
    .C(_01520_),
    .D(_01484_),
    .Y(_04549_));
 sky130_fd_sc_hd__a22o_1 _11438_ (.A1(_00454_),
    .A2(_02132_),
    .B1(_04548_),
    .B2(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__nand4_1 _11439_ (.A(_00454_),
    .B(_02132_),
    .C(_04548_),
    .D(_04549_),
    .Y(_04551_));
 sky130_fd_sc_hd__a21bo_1 _11440_ (.A1(_04038_),
    .A2(_04041_),
    .B1_N(_04039_),
    .X(_04552_));
 sky130_fd_sc_hd__and3_1 _11441_ (.A(_04550_),
    .B(_04551_),
    .C(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__a21oi_1 _11442_ (.A1(_04550_),
    .A2(_04551_),
    .B1(_04552_),
    .Y(_04554_));
 sky130_fd_sc_hd__or2_4 _11443_ (.A(_04553_),
    .B(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__or3_2 _11444_ (.A(_04047_),
    .B(_04048_),
    .C(_04050_),
    .X(_04557_));
 sky130_fd_sc_hd__nand2_1 _11445_ (.A(_00438_),
    .B(_02164_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21o_1 _11446_ (.A1(_06416_),
    .A2(_01520_),
    .B1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__xnor2_2 _11447_ (.A(_04557_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__xnor2_4 _11448_ (.A(_04555_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__or2b_1 _11449_ (.A(_04053_),
    .B_N(_04052_),
    .X(_04562_));
 sky130_fd_sc_hd__a21boi_4 _11450_ (.A1(_04046_),
    .A2(_04054_),
    .B1_N(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__xor2_4 _11451_ (.A(_04561_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__xnor2_4 _11452_ (.A(_04547_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand3_1 _11453_ (.A(_04060_),
    .B(_04078_),
    .C(_04079_),
    .Y(_04566_));
 sky130_fd_sc_hd__and2_1 _11454_ (.A(_04076_),
    .B(_04078_),
    .X(_04568_));
 sky130_fd_sc_hd__a21o_1 _11455_ (.A1(_04115_),
    .A2(_04120_),
    .B1(_04114_),
    .X(_04569_));
 sky130_fd_sc_hd__nand2_1 _11456_ (.A(_04071_),
    .B(_04075_),
    .Y(_04570_));
 sky130_fd_sc_hd__a22o_1 _11457_ (.A1(_00953_),
    .A2(net145),
    .B1(_02215_),
    .B2(_00453_),
    .X(_04571_));
 sky130_fd_sc_hd__nand4_2 _11458_ (.A(_00453_),
    .B(_00953_),
    .C(_01563_),
    .D(_02215_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand4_2 _11459_ (.A(_00985_),
    .B(_01524_),
    .C(_04571_),
    .D(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__a22o_1 _11460_ (.A1(_00985_),
    .A2(_01524_),
    .B1(_04571_),
    .B2(_04572_),
    .X(_04574_));
 sky130_fd_sc_hd__a21bo_1 _11461_ (.A1(_04065_),
    .A2(_04067_),
    .B1_N(_04066_),
    .X(_04575_));
 sky130_fd_sc_hd__a21o_1 _11462_ (.A1(_04573_),
    .A2(_04574_),
    .B1(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__nand3_1 _11463_ (.A(_04573_),
    .B(_04574_),
    .C(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__a22o_1 _11464_ (.A1(_00479_),
    .A2(_03499_),
    .B1(_04576_),
    .B2(_04577_),
    .X(_04579_));
 sky130_fd_sc_hd__nand4_1 _11465_ (.A(_00479_),
    .B(_03499_),
    .C(_04576_),
    .D(_04577_),
    .Y(_04580_));
 sky130_fd_sc_hd__a21o_1 _11466_ (.A1(_05202_),
    .A2(_01563_),
    .B1(_03532_),
    .X(_04581_));
 sky130_fd_sc_hd__and3_1 _11467_ (.A(_00062_),
    .B(_02215_),
    .C(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__nand3_1 _11468_ (.A(_04579_),
    .B(_04580_),
    .C(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__a21o_1 _11469_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__nand3_1 _11470_ (.A(_04570_),
    .B(_04583_),
    .C(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21o_1 _11471_ (.A1(_04583_),
    .A2(_04584_),
    .B1(_04570_),
    .X(_04586_));
 sky130_fd_sc_hd__and3_1 _11472_ (.A(_04569_),
    .B(_04585_),
    .C(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__a21oi_1 _11473_ (.A1(_04585_),
    .A2(_04586_),
    .B1(_04569_),
    .Y(_04588_));
 sky130_fd_sc_hd__nor3_1 _11474_ (.A(_04568_),
    .B(_04587_),
    .C(_04588_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21a_1 _11475_ (.A1(_04587_),
    .A2(_04588_),
    .B1(_04568_),
    .X(_04591_));
 sky130_fd_sc_hd__a211oi_2 _11476_ (.A1(_04566_),
    .A2(_04082_),
    .B1(_04590_),
    .C1(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__o211a_1 _11477_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04566_),
    .C1(_04082_),
    .X(_04593_));
 sky130_fd_sc_hd__nor3_2 _11478_ (.A(_04565_),
    .B(_04592_),
    .C(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__o21a_1 _11479_ (.A1(_04592_),
    .A2(_04593_),
    .B1(_04565_),
    .X(_04595_));
 sky130_fd_sc_hd__a211oi_2 _11480_ (.A1(_04533_),
    .A2(_04535_),
    .B1(_04594_),
    .C1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__o211ai_2 _11481_ (.A1(_04594_),
    .A2(_04595_),
    .B1(_04533_),
    .C1(_04535_),
    .Y(_04597_));
 sky130_fd_sc_hd__and2b_1 _11482_ (.A_N(_04596_),
    .B(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__xnor2_4 _11483_ (.A(_04532_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__and2_1 _11484_ (.A(_04130_),
    .B(_04132_),
    .X(_04601_));
 sky130_fd_sc_hd__or2_1 _11485_ (.A(_04130_),
    .B(_04132_),
    .X(_04602_));
 sky130_fd_sc_hd__o21ai_4 _11486_ (.A1(_04121_),
    .A2(_04601_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__a21oi_4 _11487_ (.A1(_04138_),
    .A2(_04164_),
    .B1(_04162_),
    .Y(_04604_));
 sky130_fd_sc_hd__a22oi_1 _11488_ (.A1(_01567_),
    .A2(_01584_),
    .B1(_02239_),
    .B2(_00481_),
    .Y(_04605_));
 sky130_fd_sc_hd__and4_1 _11489_ (.A(_00481_),
    .B(_01567_),
    .C(net188),
    .D(_02239_),
    .X(_04606_));
 sky130_fd_sc_hd__nor2_1 _11490_ (.A(_04605_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21bo_1 _11491_ (.A1(_04103_),
    .A2(_04104_),
    .B1_N(_04102_),
    .X(_04608_));
 sky130_fd_sc_hd__xor2_1 _11492_ (.A(_04607_),
    .B(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__a22oi_1 _11493_ (.A1(_01002_),
    .A2(_01562_),
    .B1(_02904_),
    .B2(_00489_),
    .Y(_04610_));
 sky130_fd_sc_hd__and4_2 _11494_ (.A(_00489_),
    .B(_01002_),
    .C(_01562_),
    .D(_02904_),
    .X(_04612_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(_04610_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__xnor2_1 _11496_ (.A(_04609_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__a21oi_1 _11497_ (.A1(_04109_),
    .A2(_04111_),
    .B1(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__and3_1 _11498_ (.A(_04109_),
    .B(_04111_),
    .C(_04614_),
    .X(_04616_));
 sky130_fd_sc_hd__nor2_2 _11499_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__xnor2_4 _11500_ (.A(_04099_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_1 _11501_ (.A(_04148_),
    .B(_04149_),
    .Y(_04619_));
 sky130_fd_sc_hd__or2b_1 _11502_ (.A(_04145_),
    .B_N(_04151_),
    .X(_04620_));
 sky130_fd_sc_hd__o21ba_1 _11503_ (.A1(_04141_),
    .A2(_04144_),
    .B1_N(_04142_),
    .X(_04621_));
 sky130_fd_sc_hd__a21oi_1 _11504_ (.A1(_04619_),
    .A2(_04620_),
    .B1(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__and3_1 _11505_ (.A(_04619_),
    .B(_04620_),
    .C(_04621_),
    .X(_04624_));
 sky130_fd_sc_hd__or2_1 _11506_ (.A(_04623_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__o21a_1 _11507_ (.A1(_03574_),
    .A2(_04124_),
    .B1(_04122_),
    .X(_04626_));
 sky130_fd_sc_hd__a21oi_1 _11508_ (.A1(_04126_),
    .A2(_04129_),
    .B1(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__nor2_1 _11509_ (.A(_04625_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__and2_1 _11510_ (.A(_04625_),
    .B(_04627_),
    .X(_04629_));
 sky130_fd_sc_hd__nor2_1 _11511_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__xnor2_2 _11512_ (.A(_04618_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__xnor2_4 _11513_ (.A(_04604_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__xor2_4 _11514_ (.A(_04603_),
    .B(_04632_),
    .X(_04634_));
 sky130_fd_sc_hd__nor2_1 _11515_ (.A(_04156_),
    .B(_04158_),
    .Y(_04635_));
 sky130_fd_sc_hd__a21o_2 _11516_ (.A1(_04152_),
    .A2(_04159_),
    .B1(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a21oi_1 _11517_ (.A1(_04167_),
    .A2(_04179_),
    .B1(_04178_),
    .Y(_04637_));
 sky130_fd_sc_hd__a22oi_1 _11518_ (.A1(_01023_),
    .A2(_01617_),
    .B1(_01603_),
    .B2(_01034_),
    .Y(_04638_));
 sky130_fd_sc_hd__and4_1 _11519_ (.A(_01034_),
    .B(_01023_),
    .C(_01617_),
    .D(_01603_),
    .X(_04639_));
 sky130_fd_sc_hd__nor2_1 _11520_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _11521_ (.A(_00507_),
    .B(_04123_),
    .Y(_04641_));
 sky130_fd_sc_hd__xor2_1 _11522_ (.A(_04640_),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_00086_),
    .B(_01617_),
    .Y(_04643_));
 sky130_fd_sc_hd__and3_1 _11524_ (.A(_00516_),
    .B(_03580_),
    .C(_04643_),
    .X(_04645_));
 sky130_fd_sc_hd__xor2_1 _11525_ (.A(_04642_),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__and3_1 _11526_ (.A(_00107_),
    .B(_04154_),
    .C(_04153_),
    .X(_04647_));
 sky130_fd_sc_hd__a31o_1 _11527_ (.A1(_00543_),
    .A2(_01629_),
    .A3(_04171_),
    .B1(_04170_),
    .X(_04648_));
 sky130_fd_sc_hd__nand2_1 _11528_ (.A(_00543_),
    .B(_04154_),
    .Y(_04649_));
 sky130_fd_sc_hd__xnor2_1 _11529_ (.A(_04648_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__xnor2_1 _11530_ (.A(_04647_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__xnor2_1 _11531_ (.A(_04646_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor2_1 _11532_ (.A(_04637_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__and2_1 _11533_ (.A(_04637_),
    .B(_04652_),
    .X(_04654_));
 sky130_fd_sc_hd__nor2_2 _11534_ (.A(_04653_),
    .B(_04654_),
    .Y(_04656_));
 sky130_fd_sc_hd__xor2_4 _11535_ (.A(_04636_),
    .B(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__a22o_1 _11536_ (.A1(_01072_),
    .A2(_01667_),
    .B1(_03019_),
    .B2(_00544_),
    .X(_04658_));
 sky130_fd_sc_hd__and4_1 _11537_ (.A(_00544_),
    .B(_01072_),
    .C(_01667_),
    .D(_03019_),
    .X(_04659_));
 sky130_fd_sc_hd__inv_2 _11538_ (.A(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__and2_1 _11539_ (.A(_04658_),
    .B(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__a21bo_1 _11540_ (.A1(_04182_),
    .A2(_04185_),
    .B1_N(_04184_),
    .X(_04662_));
 sky130_fd_sc_hd__a22oi_1 _11541_ (.A1(_01666_),
    .A2(_01652_),
    .B1(_03006_),
    .B2(_00550_),
    .Y(_04663_));
 sky130_fd_sc_hd__and4_2 _11542_ (.A(_00550_),
    .B(_01666_),
    .C(net56),
    .D(_03006_),
    .X(_04664_));
 sky130_fd_sc_hd__nor2_1 _11543_ (.A(_04663_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__xor2_1 _11544_ (.A(_04662_),
    .B(_04665_),
    .X(_04667_));
 sky130_fd_sc_hd__xor2_1 _11545_ (.A(_04193_),
    .B(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__xnor2_1 _11546_ (.A(_04661_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__a21oi_1 _11547_ (.A1(_04189_),
    .A2(_04197_),
    .B1(_04188_),
    .Y(_04670_));
 sky130_fd_sc_hd__xnor2_1 _11548_ (.A(_04669_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__and2b_1 _11549_ (.A_N(_04174_),
    .B(_04176_),
    .X(_04672_));
 sky130_fd_sc_hd__or2_2 _11550_ (.A(_03610_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__and2_1 _11551_ (.A(_04191_),
    .B(_04195_),
    .X(_04674_));
 sky130_fd_sc_hd__a21o_1 _11552_ (.A1(_03624_),
    .A2(_04196_),
    .B1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__a22o_1 _11553_ (.A1(_01051_),
    .A2(_01653_),
    .B1(net40),
    .B2(_00530_),
    .X(_04676_));
 sky130_fd_sc_hd__inv_2 _11554_ (.A(_04676_),
    .Y(_04678_));
 sky130_fd_sc_hd__and4_1 _11555_ (.A(_00530_),
    .B(_01051_),
    .C(_01653_),
    .D(_02329_),
    .X(_04679_));
 sky130_fd_sc_hd__o2bb2a_1 _11556_ (.A1_N(_01068_),
    .A2_N(_01629_),
    .B1(_04678_),
    .B2(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__and4b_1 _11557_ (.A_N(_04679_),
    .B(_01629_),
    .C(_01068_),
    .D(_04676_),
    .X(_04681_));
 sky130_fd_sc_hd__or2_1 _11558_ (.A(_04680_),
    .B(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__xnor2_1 _11559_ (.A(_04675_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__xnor2_1 _11560_ (.A(_04673_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(_04671_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__or2_1 _11562_ (.A(_04671_),
    .B(_04684_),
    .X(_04686_));
 sky130_fd_sc_hd__nand2_2 _11563_ (.A(_04685_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__and2_1 _11564_ (.A(_04198_),
    .B(_04200_),
    .X(_04689_));
 sky130_fd_sc_hd__a21oi_4 _11565_ (.A1(_04181_),
    .A2(_04201_),
    .B1(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__xor2_4 _11566_ (.A(_04687_),
    .B(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__xnor2_4 _11567_ (.A(_04657_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__or2b_1 _11568_ (.A(_04202_),
    .B_N(_04204_),
    .X(_04693_));
 sky130_fd_sc_hd__a21bo_2 _11569_ (.A1(_04165_),
    .A2(_04206_),
    .B1_N(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__xnor2_4 _11570_ (.A(_04692_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_4 _11571_ (.A(_04634_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__or2b_1 _11572_ (.A(_04207_),
    .B_N(_04209_),
    .X(_04697_));
 sky130_fd_sc_hd__a21boi_4 _11573_ (.A1(_04136_),
    .A2(_04210_),
    .B1_N(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__xnor2_4 _11574_ (.A(_04696_),
    .B(_04698_),
    .Y(_04700_));
 sky130_fd_sc_hd__xnor2_4 _11575_ (.A(_04599_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__nor2_1 _11576_ (.A(_04211_),
    .B(_04213_),
    .Y(_04702_));
 sky130_fd_sc_hd__a21oi_2 _11577_ (.A1(_04092_),
    .A2(_04214_),
    .B1(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__xor2_4 _11578_ (.A(_04701_),
    .B(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__xnor2_4 _11579_ (.A(_04531_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_1 _11580_ (.A(_04215_),
    .B(_04218_),
    .Y(_04706_));
 sky130_fd_sc_hd__a21oi_2 _11581_ (.A1(_04022_),
    .A2(_04219_),
    .B1(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__xor2_4 _11582_ (.A(_04705_),
    .B(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__xnor2_4 _11583_ (.A(_04434_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_04220_),
    .B(_04222_),
    .Y(_04711_));
 sky130_fd_sc_hd__a21oi_4 _11585_ (.A1(_03915_),
    .A2(_04223_),
    .B1(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__xor2_2 _11586_ (.A(_04709_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__xnor2_2 _11587_ (.A(_04293_),
    .B(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__nor2_1 _11588_ (.A(_04224_),
    .B(_04226_),
    .Y(_04715_));
 sky130_fd_sc_hd__a21oi_2 _11589_ (.A1(_03739_),
    .A2(_04228_),
    .B1(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__xor2_2 _11590_ (.A(_04714_),
    .B(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__xnor2_2 _11591_ (.A(_04256_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__xor2_1 _11592_ (.A(_04253_),
    .B(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__xnor2_1 _11593_ (.A(_04251_),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__and2_1 _11594_ (.A(net260),
    .B(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__nor2_1 _11595_ (.A(net260),
    .B(_04720_),
    .Y(_04722_));
 sky130_fd_sc_hd__nor2_1 _11596_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(_04243_),
    .B(_04247_),
    .Y(_04724_));
 sky130_fd_sc_hd__a21oi_1 _11598_ (.A1(_04723_),
    .A2(_04724_),
    .B1(_00166_),
    .Y(_04725_));
 sky130_fd_sc_hd__o21a_1 _11599_ (.A1(_04723_),
    .A2(_04724_),
    .B1(_04725_),
    .X(_00011_));
 sky130_fd_sc_hd__nand2_1 _11600_ (.A(net260),
    .B(_04720_),
    .Y(_04726_));
 sky130_fd_sc_hd__a31o_1 _11601_ (.A1(_04243_),
    .A2(_04247_),
    .A3(_04726_),
    .B1(_04722_),
    .X(_04727_));
 sky130_fd_sc_hd__and2b_1 _11602_ (.A_N(_04291_),
    .B(_04258_),
    .X(_04728_));
 sky130_fd_sc_hd__a21o_1 _11603_ (.A1(_04261_),
    .A2(_04290_),
    .B1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__or2b_1 _11604_ (.A(_04288_),
    .B_N(_04264_),
    .X(_04731_));
 sky130_fd_sc_hd__or2b_1 _11605_ (.A(_04263_),
    .B_N(_04289_),
    .X(_04732_));
 sky130_fd_sc_hd__and2b_1 _11606_ (.A_N(_04432_),
    .B(_04295_),
    .X(_04733_));
 sky130_fd_sc_hd__a21o_2 _11607_ (.A1(_04294_),
    .A2(_04433_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__a21o_2 _11608_ (.A1(_04265_),
    .A2(_04287_),
    .B1(_04285_),
    .X(_04735_));
 sky130_fd_sc_hd__o21ai_4 _11609_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04377_),
    .Y(_04736_));
 sky130_fd_sc_hd__a31oi_4 _11610_ (.A1(_00270_),
    .A2(_01754_),
    .A3(_04282_),
    .B1(_04279_),
    .Y(_04737_));
 sky130_fd_sc_hd__and2_1 _11611_ (.A(_04299_),
    .B(_04317_),
    .X(_04738_));
 sky130_fd_sc_hd__and2_1 _11612_ (.A(_04298_),
    .B(_04318_),
    .X(_04739_));
 sky130_fd_sc_hd__and3b_1 _11613_ (.A_N(_03709_),
    .B(_02464_),
    .C(_00617_),
    .X(_04740_));
 sky130_fd_sc_hd__xor2_1 _11614_ (.A(_04273_),
    .B(_04740_),
    .X(_04742_));
 sky130_fd_sc_hd__and2_1 _11615_ (.A(_01188_),
    .B(_01157_),
    .X(_04743_));
 sky130_fd_sc_hd__nor2_1 _11616_ (.A(_04742_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__and2_1 _11617_ (.A(_04742_),
    .B(_04743_),
    .X(_04745_));
 sky130_fd_sc_hd__or2_1 _11618_ (.A(_04744_),
    .B(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__and2b_1 _11619_ (.A_N(_03717_),
    .B(_04275_),
    .X(_04747_));
 sky130_fd_sc_hd__a31o_1 _11620_ (.A1(_01777_),
    .A2(_01157_),
    .A3(_04276_),
    .B1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__xnor2_2 _11621_ (.A(_04746_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__nand2_1 _11622_ (.A(_01777_),
    .B(_01754_),
    .Y(_04750_));
 sky130_fd_sc_hd__xnor2_1 _11623_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__o21ai_2 _11624_ (.A1(_04738_),
    .A2(_04739_),
    .B1(_04751_),
    .Y(_04753_));
 sky130_fd_sc_hd__or3_1 _11625_ (.A(_04738_),
    .B(_04739_),
    .C(_04751_),
    .X(_04754_));
 sky130_fd_sc_hd__nand2_2 _11626_ (.A(_04753_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__xor2_4 _11627_ (.A(_04737_),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__xnor2_4 _11628_ (.A(_04736_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__xnor2_4 _11629_ (.A(_04735_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__xnor2_1 _11630_ (.A(_04734_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__a21oi_1 _11631_ (.A1(_04731_),
    .A2(_04732_),
    .B1(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__and3_1 _11632_ (.A(_04731_),
    .B(_04732_),
    .C(_04759_),
    .X(_04761_));
 sky130_fd_sc_hd__nor2_1 _11633_ (.A(_04760_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__a31o_2 _11634_ (.A1(_04377_),
    .A2(_04378_),
    .A3(_04430_),
    .B1(_04429_),
    .X(_04764_));
 sky130_fd_sc_hd__a21o_2 _11635_ (.A1(_04437_),
    .A2(_04529_),
    .B1(_04528_),
    .X(_04765_));
 sky130_fd_sc_hd__or2b_1 _11636_ (.A(_04302_),
    .B_N(_04315_),
    .X(_04766_));
 sky130_fd_sc_hd__or2b_1 _11637_ (.A(_04301_),
    .B_N(_04316_),
    .X(_04767_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_04766_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__o21ai_2 _11639_ (.A1(_04335_),
    .A2(_04345_),
    .B1(_04343_),
    .Y(_04769_));
 sky130_fd_sc_hd__or2b_1 _11640_ (.A(_03759_),
    .B_N(_04313_),
    .X(_04770_));
 sky130_fd_sc_hd__o21ai_1 _11641_ (.A1(_03774_),
    .A2(_04312_),
    .B1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__and2b_1 _11642_ (.A_N(_04330_),
    .B(_04331_),
    .X(_04772_));
 sky130_fd_sc_hd__a21oi_2 _11643_ (.A1(_04332_),
    .A2(_04334_),
    .B1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__and2_1 _11644_ (.A(_01217_),
    .B(_01181_),
    .X(_04775_));
 sky130_fd_sc_hd__a21oi_1 _11645_ (.A1(_00647_),
    .A2(_02498_),
    .B1(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__and3_1 _11646_ (.A(_00647_),
    .B(_02498_),
    .C(_04775_),
    .X(_04777_));
 sky130_fd_sc_hd__nor2_1 _11647_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _11648_ (.A(_00706_),
    .B(_01784_),
    .Y(_04779_));
 sky130_fd_sc_hd__xnor2_1 _11649_ (.A(_04778_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__o21ai_2 _11650_ (.A1(_04306_),
    .A2(_04308_),
    .B1(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__or3_1 _11651_ (.A(_04306_),
    .B(_04308_),
    .C(_04780_),
    .X(_04782_));
 sky130_fd_sc_hd__and3_1 _11652_ (.A(_03772_),
    .B(_04781_),
    .C(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__a21oi_1 _11653_ (.A1(_04781_),
    .A2(_04782_),
    .B1(_03772_),
    .Y(_04784_));
 sky130_fd_sc_hd__or2_1 _11654_ (.A(_04783_),
    .B(_04784_),
    .X(_04786_));
 sky130_fd_sc_hd__xnor2_2 _11655_ (.A(_04310_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__xnor2_1 _11656_ (.A(_04773_),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__xnor2_1 _11657_ (.A(_04771_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__xnor2_1 _11658_ (.A(_04769_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__xor2_1 _11659_ (.A(_04768_),
    .B(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__or2b_1 _11660_ (.A(_04327_),
    .B_N(_04326_),
    .X(_04792_));
 sky130_fd_sc_hd__nand3_1 _11661_ (.A(_00200_),
    .B(_03180_),
    .C(_04328_),
    .Y(_04793_));
 sky130_fd_sc_hd__a22o_1 _11662_ (.A1(_01251_),
    .A2(_01835_),
    .B1(_01858_),
    .B2(_00703_),
    .X(_04794_));
 sky130_fd_sc_hd__nand4_1 _11663_ (.A(_00703_),
    .B(_01251_),
    .C(_01835_),
    .D(_01858_),
    .Y(_04795_));
 sky130_fd_sc_hd__a31o_1 _11664_ (.A1(_00672_),
    .A2(_01835_),
    .A3(_04320_),
    .B1(_04321_),
    .X(_04797_));
 sky130_fd_sc_hd__and3_1 _11665_ (.A(_04794_),
    .B(_04795_),
    .C(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__a21oi_1 _11666_ (.A1(_04794_),
    .A2(_04795_),
    .B1(_04797_),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_1 _11667_ (.A(_04798_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _11668_ (.A(_00672_),
    .B(_03180_),
    .Y(_04801_));
 sky130_fd_sc_hd__xor2_1 _11669_ (.A(_04800_),
    .B(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__a21oi_2 _11670_ (.A1(_04792_),
    .A2(_04793_),
    .B1(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__and3_1 _11671_ (.A(_04792_),
    .B(_04793_),
    .C(_04802_),
    .X(_04804_));
 sky130_fd_sc_hd__or2_1 _11672_ (.A(_04803_),
    .B(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__a22o_1 _11673_ (.A1(_03817_),
    .A2(_03826_),
    .B1(_04339_),
    .B2(_04341_),
    .X(_04806_));
 sky130_fd_sc_hd__nor2_1 _11674_ (.A(_04354_),
    .B(_04361_),
    .Y(_04808_));
 sky130_fd_sc_hd__and2_1 _11675_ (.A(_04354_),
    .B(_04361_),
    .X(_04809_));
 sky130_fd_sc_hd__a2bb2o_1 _11676_ (.A1_N(_04808_),
    .A2_N(_04809_),
    .B1(_04355_),
    .B2(_04363_),
    .X(_04810_));
 sky130_fd_sc_hd__xnor2_1 _11677_ (.A(_04806_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__or2_1 _11678_ (.A(_04805_),
    .B(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_04805_),
    .B(_04811_),
    .Y(_04813_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(_04812_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__and2_1 _11681_ (.A(_03881_),
    .B(_04397_),
    .X(_04815_));
 sky130_fd_sc_hd__a32o_1 _11682_ (.A1(_00291_),
    .A2(_02592_),
    .A3(_04390_),
    .B1(_04389_),
    .B2(_01309_),
    .X(_04816_));
 sky130_fd_sc_hd__and2_1 _11683_ (.A(_00201_),
    .B(_01264_),
    .X(_04817_));
 sky130_fd_sc_hd__a22oi_1 _11684_ (.A1(_01264_),
    .A2(_01250_),
    .B1(_03210_),
    .B2(_00677_),
    .Y(_04819_));
 sky130_fd_sc_hd__and4_1 _11685_ (.A(_00677_),
    .B(_01264_),
    .C(_01250_),
    .D(_03210_),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _11686_ (.A(_00665_),
    .B(_01872_),
    .Y(_04821_));
 sky130_fd_sc_hd__or4_1 _11687_ (.A(_04817_),
    .B(_04819_),
    .C(_04820_),
    .D(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__o22ai_1 _11688_ (.A1(_04819_),
    .A2(_04820_),
    .B1(_04821_),
    .B2(_04817_),
    .Y(_04823_));
 sky130_fd_sc_hd__and3_1 _11689_ (.A(_04816_),
    .B(_04822_),
    .C(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__a21oi_1 _11690_ (.A1(_04822_),
    .A2(_04823_),
    .B1(_04816_),
    .Y(_04825_));
 sky130_fd_sc_hd__nor2_1 _11691_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__o21ai_1 _11692_ (.A1(_04815_),
    .A2(_04400_),
    .B1(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__or3_1 _11693_ (.A(_04815_),
    .B(_04400_),
    .C(_04826_),
    .X(_04828_));
 sky130_fd_sc_hd__and2_1 _11694_ (.A(_04827_),
    .B(_04828_),
    .X(_04830_));
 sky130_fd_sc_hd__xnor2_2 _11695_ (.A(_04365_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__or2b_1 _11696_ (.A(_04367_),
    .B_N(_04350_),
    .X(_04832_));
 sky130_fd_sc_hd__a21bo_1 _11697_ (.A1(_04349_),
    .A2(_04368_),
    .B1_N(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__xor2_2 _11698_ (.A(_04831_),
    .B(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__xnor2_2 _11699_ (.A(_04814_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__and2b_1 _11700_ (.A_N(_04370_),
    .B(_04372_),
    .X(_04836_));
 sky130_fd_sc_hd__a21oi_2 _11701_ (.A1(_04346_),
    .A2(_04373_),
    .B1(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__xnor2_1 _11702_ (.A(_04835_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nor2_1 _11703_ (.A(_04791_),
    .B(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__and2_1 _11704_ (.A(_04791_),
    .B(_04838_),
    .X(_04841_));
 sky130_fd_sc_hd__nor2_4 _11705_ (.A(_04839_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__and2b_1 _11706_ (.A_N(_04422_),
    .B(_04386_),
    .X(_04843_));
 sky130_fd_sc_hd__a21o_2 _11707_ (.A1(_04388_),
    .A2(_04421_),
    .B1(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__or2b_1 _11708_ (.A(_04486_),
    .B_N(_04488_),
    .X(_04845_));
 sky130_fd_sc_hd__a21boi_2 _11709_ (.A1(_04455_),
    .A2(_04489_),
    .B1_N(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__or2b_1 _11710_ (.A(_04417_),
    .B_N(_04419_),
    .X(_04847_));
 sky130_fd_sc_hd__a21bo_2 _11711_ (.A1(_04403_),
    .A2(_04420_),
    .B1_N(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__nor2_1 _11712_ (.A(_04441_),
    .B(_04453_),
    .Y(_04849_));
 sky130_fd_sc_hd__a21o_1 _11713_ (.A1(_04440_),
    .A2(_04454_),
    .B1(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__inv_2 _11714_ (.A(_03868_),
    .Y(_04852_));
 sky130_fd_sc_hd__and2b_1 _11715_ (.A_N(_04394_),
    .B(_04396_),
    .X(_04853_));
 sky130_fd_sc_hd__and3_1 _11716_ (.A(_00343_),
    .B(_03859_),
    .C(_04404_),
    .X(_04854_));
 sky130_fd_sc_hd__a22o_1 _11717_ (.A1(_01309_),
    .A2(_01288_),
    .B1(_02615_),
    .B2(_00749_),
    .X(_04855_));
 sky130_fd_sc_hd__nand4_2 _11718_ (.A(_00749_),
    .B(_01309_),
    .C(_01288_),
    .D(_02615_),
    .Y(_04856_));
 sky130_fd_sc_hd__a22o_1 _11719_ (.A1(_00774_),
    .A2(_02592_),
    .B1(_04855_),
    .B2(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__nand4_2 _11720_ (.A(_00774_),
    .B(_02592_),
    .C(_04855_),
    .D(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _11721_ (.A(_04857_),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__xnor2_1 _11722_ (.A(_04854_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__o21a_1 _11723_ (.A1(_04852_),
    .A2(_04853_),
    .B1(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__nor3_1 _11724_ (.A(_04852_),
    .B(_04853_),
    .C(_04860_),
    .Y(_04863_));
 sky130_fd_sc_hd__or2_2 _11725_ (.A(_04861_),
    .B(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__a22o_1 _11726_ (.A1(_01365_),
    .A2(_02626_),
    .B1(_01986_),
    .B2(_00757_),
    .X(_04865_));
 sky130_fd_sc_hd__nand4_1 _11727_ (.A(_00757_),
    .B(_01365_),
    .C(_02626_),
    .D(_01986_),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_2 _11728_ (.A(_04865_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__and3_1 _11729_ (.A(_00810_),
    .B(_02626_),
    .C(_04409_),
    .X(_04868_));
 sky130_fd_sc_hd__o211a_2 _11730_ (.A1(_04408_),
    .A2(_04868_),
    .B1(_00810_),
    .C1(_03859_),
    .X(_04869_));
 sky130_fd_sc_hd__a211oi_1 _11731_ (.A1(_00810_),
    .A2(_03859_),
    .B1(_04408_),
    .C1(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_2 _11732_ (.A(_04869_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__xor2_4 _11733_ (.A(_04867_),
    .B(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__a21o_2 _11734_ (.A1(_04411_),
    .A2(_04412_),
    .B1(_04415_),
    .X(_04874_));
 sky130_fd_sc_hd__xor2_4 _11735_ (.A(_04872_),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__xor2_4 _11736_ (.A(_04864_),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__xor2_2 _11737_ (.A(_04850_),
    .B(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__xnor2_2 _11738_ (.A(_04848_),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__xor2_2 _11739_ (.A(_04846_),
    .B(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__xnor2_1 _11740_ (.A(_04844_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _11741_ (.A(_04384_),
    .B(_04423_),
    .Y(_04881_));
 sky130_fd_sc_hd__a21oi_2 _11742_ (.A1(_04382_),
    .A2(_04425_),
    .B1(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nor2_1 _11743_ (.A(_04880_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__and2_1 _11744_ (.A(_04880_),
    .B(_04882_),
    .X(_04885_));
 sky130_fd_sc_hd__nor2_2 _11745_ (.A(_04883_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__xor2_4 _11746_ (.A(_04842_),
    .B(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__xor2_4 _11747_ (.A(_04765_),
    .B(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__xor2_4 _11748_ (.A(_04764_),
    .B(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__nor2_1 _11749_ (.A(_04522_),
    .B(_04525_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21o_1 _11750_ (.A1(_04491_),
    .A2(_04526_),
    .B1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__a21oi_2 _11751_ (.A1(_04532_),
    .A2(_04597_),
    .B1(_04596_),
    .Y(_04892_));
 sky130_fd_sc_hd__and3_1 _11752_ (.A(_04448_),
    .B(_04449_),
    .C(_04452_),
    .X(_04893_));
 sky130_fd_sc_hd__a21oi_1 _11753_ (.A1(_04459_),
    .A2(_04472_),
    .B1(_04471_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand2_1 _11754_ (.A(_01385_),
    .B(_01987_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _11755_ (.A(_02694_),
    .B(_01367_),
    .Y(_04897_));
 sky130_fd_sc_hd__xor2_1 _11756_ (.A(_04896_),
    .B(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__xor2_1 _11757_ (.A(_04458_),
    .B(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__xnor2_1 _11758_ (.A(_04443_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__a21oi_1 _11759_ (.A1(_04445_),
    .A2(_04449_),
    .B1(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__and3_1 _11760_ (.A(_04445_),
    .B(_04449_),
    .C(_04900_),
    .X(_04902_));
 sky130_fd_sc_hd__or2_1 _11761_ (.A(_04901_),
    .B(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__xor2_1 _11762_ (.A(_04894_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nor2_1 _11763_ (.A(_04893_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__and2_1 _11764_ (.A(_04893_),
    .B(_04904_),
    .X(_04907_));
 sky130_fd_sc_hd__or2_1 _11765_ (.A(_04905_),
    .B(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__and2_1 _11766_ (.A(_00830_),
    .B(_02695_),
    .X(_04909_));
 sky130_fd_sc_hd__and4_1 _11767_ (.A(_00821_),
    .B(_01410_),
    .C(_01397_),
    .D(_02731_),
    .X(_04910_));
 sky130_fd_sc_hd__a22oi_2 _11768_ (.A1(_01410_),
    .A2(_01397_),
    .B1(_02731_),
    .B2(_00821_),
    .Y(_04911_));
 sky130_fd_sc_hd__nor2_1 _11769_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__nand2_1 _11770_ (.A(_00850_),
    .B(_02019_),
    .Y(_04913_));
 sky130_fd_sc_hd__xnor2_1 _11771_ (.A(_04912_),
    .B(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__and2_1 _11772_ (.A(_04461_),
    .B(_04463_),
    .X(_04915_));
 sky130_fd_sc_hd__xor2_1 _11773_ (.A(_04914_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__a21bo_1 _11774_ (.A1(_04465_),
    .A2(_04466_),
    .B1_N(_04464_),
    .X(_04918_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(_04916_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__nor2_1 _11776_ (.A(_04909_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__and2_1 _11777_ (.A(_04909_),
    .B(_04919_),
    .X(_04921_));
 sky130_fd_sc_hd__or2_1 _11778_ (.A(_04920_),
    .B(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__and2_1 _11779_ (.A(_04505_),
    .B(_04506_),
    .X(_04923_));
 sky130_fd_sc_hd__nand2_1 _11780_ (.A(_00879_),
    .B(_03967_),
    .Y(_04924_));
 sky130_fd_sc_hd__xnor2_1 _11781_ (.A(_04923_),
    .B(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__nor2_1 _11782_ (.A(_04476_),
    .B(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__and2_1 _11783_ (.A(_04476_),
    .B(_04925_),
    .X(_04927_));
 sky130_fd_sc_hd__or2_2 _11784_ (.A(_04926_),
    .B(_04927_),
    .X(_04929_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_03966_),
    .B(_04480_),
    .Y(_04930_));
 sky130_fd_sc_hd__o31a_1 _11786_ (.A1(_04475_),
    .A2(_04476_),
    .A3(_04477_),
    .B1(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__xnor2_2 _11787_ (.A(_04929_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__xnor2_2 _11788_ (.A(_04922_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _11789_ (.A(_04481_),
    .B(_04484_),
    .Y(_04934_));
 sky130_fd_sc_hd__o21a_1 _11790_ (.A1(_04474_),
    .A2(_04485_),
    .B1(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__xnor2_2 _11791_ (.A(_04933_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__xor2_1 _11792_ (.A(_04908_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_04499_),
    .B(_04518_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21bo_2 _11794_ (.A1(_04497_),
    .A2(_04519_),
    .B1_N(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_1 _11795_ (.A(_04561_),
    .B(_04563_),
    .Y(_04941_));
 sky130_fd_sc_hd__a21o_1 _11796_ (.A1(_04547_),
    .A2(_04564_),
    .B1(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__nor2_1 _11797_ (.A(_04507_),
    .B(_04517_),
    .Y(_04943_));
 sky130_fd_sc_hd__a21o_2 _11798_ (.A1(_04508_),
    .A2(_04516_),
    .B1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__nor2_1 _11799_ (.A(_04044_),
    .B(_04045_),
    .Y(_04945_));
 sky130_fd_sc_hd__a21o_1 _11800_ (.A1(_04945_),
    .A2(_04542_),
    .B1(_04546_),
    .X(_04946_));
 sky130_fd_sc_hd__a22oi_1 _11801_ (.A1(_01444_),
    .A2(_01434_),
    .B1(_02765_),
    .B2(_00872_),
    .Y(_04947_));
 sky130_fd_sc_hd__and4_1 _11802_ (.A(_00872_),
    .B(_01444_),
    .C(_01434_),
    .D(_02765_),
    .X(_04948_));
 sky130_fd_sc_hd__or2_2 _11803_ (.A(_04947_),
    .B(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__a32o_2 _11804_ (.A1(_00879_),
    .A2(_01434_),
    .A3(_04502_),
    .B1(_04500_),
    .B2(_02765_),
    .X(_04951_));
 sky130_fd_sc_hd__xnor2_4 _11805_ (.A(_04949_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__and2_1 _11806_ (.A(_01488_),
    .B(_01443_),
    .X(_04953_));
 sky130_fd_sc_hd__and3_1 _11807_ (.A(_01487_),
    .B(_02064_),
    .C(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__nand2_1 _11808_ (.A(_04511_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(_04511_),
    .B(_04954_),
    .X(_04956_));
 sky130_fd_sc_hd__a21o_1 _11810_ (.A1(_01487_),
    .A2(_02064_),
    .B1(_04953_),
    .X(_04957_));
 sky130_fd_sc_hd__and3_1 _11811_ (.A(_04955_),
    .B(_04956_),
    .C(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__xnor2_2 _11812_ (.A(_04515_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__xnor2_4 _11813_ (.A(_04952_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__xnor2_2 _11814_ (.A(_04946_),
    .B(_04960_),
    .Y(_04962_));
 sky130_fd_sc_hd__xor2_2 _11815_ (.A(_04944_),
    .B(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__xor2_2 _11816_ (.A(_04942_),
    .B(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__xor2_4 _11817_ (.A(_04940_),
    .B(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__and2b_1 _11818_ (.A_N(_04520_),
    .B(_04495_),
    .X(_04966_));
 sky130_fd_sc_hd__a21o_1 _11819_ (.A1(_04493_),
    .A2(_04521_),
    .B1(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__xor2_1 _11820_ (.A(_04965_),
    .B(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__xnor2_1 _11821_ (.A(_04937_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__xor2_1 _11822_ (.A(_04892_),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__nand2_1 _11823_ (.A(_04891_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__or2_1 _11824_ (.A(_04891_),
    .B(_04970_),
    .X(_04973_));
 sky130_fd_sc_hd__and2_2 _11825_ (.A(_04971_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__or2_1 _11826_ (.A(_04592_),
    .B(_04594_),
    .X(_04975_));
 sky130_fd_sc_hd__or2b_1 _11827_ (.A(_04604_),
    .B_N(_04631_),
    .X(_04976_));
 sky130_fd_sc_hd__a21boi_4 _11828_ (.A1(_04603_),
    .A2(_04632_),
    .B1_N(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__or2b_1 _11829_ (.A(_04540_),
    .B_N(_04541_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_1 _11830_ (.A(_00421_),
    .B(_01488_),
    .Y(_04979_));
 sky130_fd_sc_hd__and3_1 _11831_ (.A(_00937_),
    .B(_02799_),
    .C(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__xnor2_1 _11832_ (.A(_04553_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _11833_ (.A(_04978_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__or2_1 _11834_ (.A(_04978_),
    .B(_04981_),
    .X(_04984_));
 sky130_fd_sc_hd__nand2_2 _11835_ (.A(_04982_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__a22o_1 _11836_ (.A1(_01520_),
    .A2(_01484_),
    .B1(_02164_),
    .B2(_00910_),
    .X(_04986_));
 sky130_fd_sc_hd__nand4_1 _11837_ (.A(_00910_),
    .B(_01520_),
    .C(_01484_),
    .D(_02164_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _11838_ (.A(_04986_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _11839_ (.A(_00956_),
    .B(_02132_),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_1 _11840_ (.A(_04988_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _11841_ (.A(_04549_),
    .B(_04551_),
    .Y(_04991_));
 sky130_fd_sc_hd__xnor2_1 _11842_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_1 _11843_ (.A(_04048_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__or2_1 _11844_ (.A(_04048_),
    .B(_04992_),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_2 _11845_ (.A(_04993_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__and2_1 _11846_ (.A(_04557_),
    .B(_04559_),
    .X(_04997_));
 sky130_fd_sc_hd__or2_1 _11847_ (.A(_04557_),
    .B(_04559_),
    .X(_04998_));
 sky130_fd_sc_hd__o21ai_4 _11848_ (.A1(_04555_),
    .A2(_04997_),
    .B1(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__xor2_4 _11849_ (.A(_04996_),
    .B(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__xor2_4 _11850_ (.A(_04985_),
    .B(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__o21ba_1 _11851_ (.A1(_04568_),
    .A2(_04588_),
    .B1_N(_04587_),
    .X(_05002_));
 sky130_fd_sc_hd__nand2_1 _11852_ (.A(_04583_),
    .B(_04585_),
    .Y(_05003_));
 sky130_fd_sc_hd__a21o_1 _11853_ (.A1(_04109_),
    .A2(_04111_),
    .B1(_04614_),
    .X(_05004_));
 sky130_fd_sc_hd__o21ai_2 _11854_ (.A1(_04100_),
    .A2(_04616_),
    .B1(_05004_),
    .Y(_05006_));
 sky130_fd_sc_hd__a22o_1 _11855_ (.A1(_01563_),
    .A2(_01524_),
    .B1(_02215_),
    .B2(_00953_),
    .X(_05007_));
 sky130_fd_sc_hd__nand4_1 _11856_ (.A(_00953_),
    .B(_01563_),
    .C(_01524_),
    .D(_02215_),
    .Y(_05008_));
 sky130_fd_sc_hd__nand2_1 _11857_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_1 _11858_ (.A(_04572_),
    .B(_04573_),
    .Y(_05010_));
 sky130_fd_sc_hd__xnor2_2 _11859_ (.A(_05009_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _11860_ (.A(_00985_),
    .B(_03499_),
    .Y(_05012_));
 sky130_fd_sc_hd__xor2_2 _11861_ (.A(_05011_),
    .B(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__and2_1 _11862_ (.A(_04577_),
    .B(_04580_),
    .X(_05014_));
 sky130_fd_sc_hd__xnor2_1 _11863_ (.A(_05013_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__xnor2_1 _11864_ (.A(_05006_),
    .B(_05015_),
    .Y(_05017_));
 sky130_fd_sc_hd__xor2_1 _11865_ (.A(_05003_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__and2b_1 _11866_ (.A_N(_05002_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__and2b_1 _11867_ (.A_N(_05018_),
    .B(_05002_),
    .X(_05020_));
 sky130_fd_sc_hd__nor2_1 _11868_ (.A(_05019_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__xnor2_2 _11869_ (.A(_05001_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__xor2_2 _11870_ (.A(_04977_),
    .B(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__xor2_2 _11871_ (.A(_04975_),
    .B(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__or2_1 _11872_ (.A(_04625_),
    .B(_04627_),
    .X(_05025_));
 sky130_fd_sc_hd__o21ai_4 _11873_ (.A1(_04618_),
    .A2(_04629_),
    .B1(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__a21o_2 _11874_ (.A1(_04636_),
    .A2(_04656_),
    .B1(_04653_),
    .X(_05028_));
 sky130_fd_sc_hd__nand2_1 _11875_ (.A(_04607_),
    .B(_04608_),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _11876_ (.A(_04609_),
    .B(_04613_),
    .Y(_05030_));
 sky130_fd_sc_hd__a22oi_1 _11877_ (.A1(_01584_),
    .A2(_01562_),
    .B1(_02904_),
    .B2(_01002_),
    .Y(_05031_));
 sky130_fd_sc_hd__and4_1 _11878_ (.A(_01002_),
    .B(_01584_),
    .C(_01562_),
    .D(_02904_),
    .X(_05032_));
 sky130_fd_sc_hd__nor2_1 _11879_ (.A(_05031_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(_00481_),
    .B(_01584_),
    .Y(_05034_));
 sky130_fd_sc_hd__and3_1 _11881_ (.A(_01567_),
    .B(_02239_),
    .C(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__xnor2_1 _11882_ (.A(_05033_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__a21o_1 _11883_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__nand3_1 _11884_ (.A(_05029_),
    .B(_05030_),
    .C(_05036_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_2 _11885_ (.A(_05037_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__xor2_4 _11886_ (.A(_04612_),
    .B(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__and2b_1 _11887_ (.A_N(_04642_),
    .B(_04645_),
    .X(_05042_));
 sky130_fd_sc_hd__or2_1 _11888_ (.A(_04147_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__and3_1 _11889_ (.A(_00507_),
    .B(_04123_),
    .C(_04640_),
    .X(_05044_));
 sky130_fd_sc_hd__nor2_1 _11890_ (.A(_04639_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__xnor2_1 _11891_ (.A(_05043_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2_1 _11892_ (.A(_04623_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__or2_1 _11893_ (.A(_04623_),
    .B(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_2 _11894_ (.A(_05047_),
    .B(_05048_),
    .Y(_05050_));
 sky130_fd_sc_hd__xor2_4 _11895_ (.A(_05041_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__xor2_4 _11896_ (.A(_05028_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__xnor2_4 _11897_ (.A(_05026_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__and2_2 _11898_ (.A(_04661_),
    .B(_04668_),
    .X(_05054_));
 sky130_fd_sc_hd__nand2_2 _11899_ (.A(_01072_),
    .B(_03019_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_2 _11900_ (.A(_01666_),
    .B(_03006_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_2 _11901_ (.A(_01667_),
    .B(_01652_),
    .Y(_05057_));
 sky130_fd_sc_hd__xor2_4 _11902_ (.A(_05056_),
    .B(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__xnor2_4 _11903_ (.A(_04660_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__xor2_4 _11904_ (.A(_04664_),
    .B(_05059_),
    .X(_05061_));
 sky130_fd_sc_hd__xnor2_4 _11905_ (.A(_05055_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__xnor2_4 _11906_ (.A(_05054_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _11907_ (.A(_04662_),
    .B(_04665_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand2_1 _11908_ (.A(_04193_),
    .B(_04667_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand2_2 _11909_ (.A(_05064_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__a22oi_1 _11910_ (.A1(_01653_),
    .A2(_01629_),
    .B1(_02329_),
    .B2(_01051_),
    .Y(_05067_));
 sky130_fd_sc_hd__and4_1 _11911_ (.A(_01051_),
    .B(_01653_),
    .C(_01629_),
    .D(_02329_),
    .X(_05068_));
 sky130_fd_sc_hd__nor2_2 _11912_ (.A(_05067_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__xor2_4 _11913_ (.A(_05066_),
    .B(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__xnor2_4 _11914_ (.A(_05063_),
    .B(_05070_),
    .Y(_05072_));
 sky130_fd_sc_hd__o21a_2 _11915_ (.A1(_04669_),
    .A2(_04670_),
    .B1(_04686_),
    .X(_05073_));
 sky130_fd_sc_hd__xnor2_4 _11916_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_04647_),
    .B(_04650_),
    .Y(_05075_));
 sky130_fd_sc_hd__o21ai_1 _11918_ (.A1(_04646_),
    .A2(_04651_),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__or2b_1 _11919_ (.A(_04682_),
    .B_N(_04675_),
    .X(_05077_));
 sky130_fd_sc_hd__a21bo_1 _11920_ (.A1(_04673_),
    .A2(_04683_),
    .B1_N(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a22o_1 _11921_ (.A1(_01617_),
    .A2(_01603_),
    .B1(_03580_),
    .B2(_01023_),
    .X(_05079_));
 sky130_fd_sc_hd__nand4_2 _11922_ (.A(_01023_),
    .B(_01617_),
    .C(_01603_),
    .D(_03580_),
    .Y(_05080_));
 sky130_fd_sc_hd__a22o_1 _11923_ (.A1(_01034_),
    .A2(_04123_),
    .B1(_05079_),
    .B2(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__nand4_1 _11924_ (.A(_01034_),
    .B(_04123_),
    .C(_05079_),
    .D(_05080_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _11925_ (.A(_05081_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__and3_1 _11926_ (.A(_00543_),
    .B(_04154_),
    .C(_04648_),
    .X(_05085_));
 sky130_fd_sc_hd__nor2_1 _11927_ (.A(_04679_),
    .B(_04681_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_2 _11928_ (.A(_01068_),
    .B(_04154_),
    .Y(_05087_));
 sky130_fd_sc_hd__xnor2_1 _11929_ (.A(_05086_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__xor2_1 _11930_ (.A(_05085_),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__xor2_1 _11931_ (.A(_05084_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__xor2_1 _11932_ (.A(_05078_),
    .B(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__and2_1 _11933_ (.A(_05076_),
    .B(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__nor2_1 _11934_ (.A(_05076_),
    .B(_05091_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_2 _11935_ (.A(_05092_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__xnor2_4 _11936_ (.A(_05074_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nor2_1 _11937_ (.A(_04687_),
    .B(_04690_),
    .Y(_05097_));
 sky130_fd_sc_hd__a21oi_4 _11938_ (.A1(_04657_),
    .A2(_04691_),
    .B1(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__xnor2_4 _11939_ (.A(_05096_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_4 _11940_ (.A(_05053_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__or2b_1 _11941_ (.A(_04692_),
    .B_N(_04694_),
    .X(_05101_));
 sky130_fd_sc_hd__a21boi_4 _11942_ (.A1(_04634_),
    .A2(_04695_),
    .B1_N(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xor2_2 _11943_ (.A(_05100_),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__xnor2_2 _11944_ (.A(_05024_),
    .B(_05103_),
    .Y(_05105_));
 sky130_fd_sc_hd__or2_1 _11945_ (.A(_04696_),
    .B(_04698_),
    .X(_05106_));
 sky130_fd_sc_hd__o21a_2 _11946_ (.A1(_04599_),
    .A2(_04700_),
    .B1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__xor2_2 _11947_ (.A(_05105_),
    .B(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__xnor2_2 _11948_ (.A(_04974_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__nor2_1 _11949_ (.A(_04701_),
    .B(_04703_),
    .Y(_05110_));
 sky130_fd_sc_hd__a21oi_2 _11950_ (.A1(_04531_),
    .A2(_04704_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__xor2_2 _11951_ (.A(_05109_),
    .B(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__xnor2_2 _11952_ (.A(_04889_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_04705_),
    .B(_04707_),
    .Y(_05114_));
 sky130_fd_sc_hd__a21oi_2 _11954_ (.A1(_04434_),
    .A2(_04708_),
    .B1(_05114_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _11955_ (.A(_05113_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_05113_),
    .B(_05116_),
    .Y(_05118_));
 sky130_fd_sc_hd__and2b_1 _11957_ (.A_N(_05117_),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__xnor2_1 _11958_ (.A(_04762_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__nor2_1 _11959_ (.A(_04709_),
    .B(_04712_),
    .Y(_05121_));
 sky130_fd_sc_hd__a21oi_1 _11960_ (.A1(_04293_),
    .A2(_04713_),
    .B1(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__xnor2_1 _11961_ (.A(_05120_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__xor2_1 _11962_ (.A(_04729_),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__nor2_1 _11963_ (.A(_04714_),
    .B(_04716_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_1 _11964_ (.A1(_04256_),
    .A2(_04717_),
    .B1(_05125_),
    .Y(_05127_));
 sky130_fd_sc_hd__or2_1 _11965_ (.A(_05124_),
    .B(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_05124_),
    .B(_05127_),
    .Y(_05129_));
 sky130_fd_sc_hd__and2_1 _11967_ (.A(_05128_),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__and2_1 _11968_ (.A(_04236_),
    .B(_04719_),
    .X(_05131_));
 sky130_fd_sc_hd__nand2_1 _11969_ (.A(_04253_),
    .B(_04718_),
    .Y(_05132_));
 sky130_fd_sc_hd__nor2_1 _11970_ (.A(_04253_),
    .B(_04718_),
    .Y(_05133_));
 sky130_fd_sc_hd__a221o_1 _11971_ (.A1(_04250_),
    .A2(_05132_),
    .B1(_05131_),
    .B2(_04240_),
    .C1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__a31o_4 _11972_ (.A1(_03065_),
    .A2(_04237_),
    .A3(_05131_),
    .B1(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__xor2_1 _11973_ (.A(_05130_),
    .B(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(net261),
    .B(_05136_),
    .Y(_05138_));
 sky130_fd_sc_hd__or2_1 _11975_ (.A(net261),
    .B(_05136_),
    .X(_05139_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_05138_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(_04727_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__or2_1 _11978_ (.A(_04727_),
    .B(_05140_),
    .X(_05142_));
 sky130_fd_sc_hd__and3_1 _11979_ (.A(_02185_),
    .B(_05141_),
    .C(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_1 _11980_ (.A(_05143_),
    .X(_00012_));
 sky130_fd_sc_hd__a21boi_2 _11981_ (.A1(_05130_),
    .A2(_05135_),
    .B1_N(_05128_),
    .Y(_05144_));
 sky130_fd_sc_hd__or2_1 _11982_ (.A(_05120_),
    .B(_05122_),
    .X(_05145_));
 sky130_fd_sc_hd__or2b_1 _11983_ (.A(_05123_),
    .B_N(_04729_),
    .X(_05146_));
 sky130_fd_sc_hd__a21o_1 _11984_ (.A1(_04734_),
    .A2(_04758_),
    .B1(_04760_),
    .X(_05148_));
 sky130_fd_sc_hd__and2_1 _11985_ (.A(_04765_),
    .B(_04887_),
    .X(_05149_));
 sky130_fd_sc_hd__a21o_1 _11986_ (.A1(_04764_),
    .A2(_04888_),
    .B1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__o21ai_4 _11987_ (.A1(_04737_),
    .A2(_04755_),
    .B1(_04753_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21bai_4 _11988_ (.A1(_04835_),
    .A2(_04837_),
    .B1_N(_04839_),
    .Y(_05152_));
 sky130_fd_sc_hd__and2b_1 _11989_ (.A_N(_04746_),
    .B(_04748_),
    .X(_05153_));
 sky130_fd_sc_hd__a31oi_4 _11990_ (.A1(_01777_),
    .A2(_01754_),
    .A3(_04749_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_1 _11991_ (.A(_04769_),
    .B(_04789_),
    .Y(_05155_));
 sky130_fd_sc_hd__or2b_1 _11992_ (.A(_04790_),
    .B_N(_04768_),
    .X(_05156_));
 sky130_fd_sc_hd__a21o_1 _11993_ (.A1(_04273_),
    .A2(_04740_),
    .B1(_04745_),
    .X(_05157_));
 sky130_fd_sc_hd__and3_1 _11994_ (.A(_00617_),
    .B(_02464_),
    .C(_03709_),
    .X(_05159_));
 sky130_fd_sc_hd__nand2_1 _11995_ (.A(_01157_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a21o_1 _11996_ (.A1(_01157_),
    .A2(_02464_),
    .B1(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_05160_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__xnor2_1 _11998_ (.A(_05157_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_1 _11999_ (.A(_01188_),
    .B(_01754_),
    .Y(_05164_));
 sky130_fd_sc_hd__xor2_1 _12000_ (.A(_05163_),
    .B(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__a21o_1 _12001_ (.A1(_05155_),
    .A2(_05156_),
    .B1(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__nand3_1 _12002_ (.A(_05155_),
    .B(_05156_),
    .C(_05165_),
    .Y(_05167_));
 sky130_fd_sc_hd__and2_1 _12003_ (.A(_05166_),
    .B(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__xnor2_2 _12004_ (.A(_05154_),
    .B(_05168_),
    .Y(_05170_));
 sky130_fd_sc_hd__xnor2_2 _12005_ (.A(_05152_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__xnor2_4 _12006_ (.A(_05151_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__xnor2_1 _12007_ (.A(_05150_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__and2b_1 _12008_ (.A_N(_04757_),
    .B(_04735_),
    .X(_05174_));
 sky130_fd_sc_hd__a21o_2 _12009_ (.A1(_04736_),
    .A2(_04756_),
    .B1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__and2b_1 _12010_ (.A_N(_05173_),
    .B(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__and2b_1 _12011_ (.A_N(_05175_),
    .B(_05173_),
    .X(_05177_));
 sky130_fd_sc_hd__nor2_1 _12012_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a21o_1 _12013_ (.A1(_04842_),
    .A2(_04886_),
    .B1(_04883_),
    .X(_05179_));
 sky130_fd_sc_hd__o21a_1 _12014_ (.A1(_04892_),
    .A2(_04969_),
    .B1(_04971_),
    .X(_05181_));
 sky130_fd_sc_hd__or2b_1 _12015_ (.A(_04788_),
    .B_N(_04771_),
    .X(_05182_));
 sky130_fd_sc_hd__o21ai_4 _12016_ (.A1(_04773_),
    .A2(_04787_),
    .B1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21bo_2 _12017_ (.A1(_04806_),
    .A2(_04810_),
    .B1_N(_04812_),
    .X(_05184_));
 sky130_fd_sc_hd__nor2_1 _12018_ (.A(_04310_),
    .B(_04786_),
    .Y(_05185_));
 sky130_fd_sc_hd__a22oi_1 _12019_ (.A1(_01181_),
    .A2(_02498_),
    .B1(_01784_),
    .B2(_01217_),
    .Y(_05186_));
 sky130_fd_sc_hd__a31o_1 _12020_ (.A1(_02498_),
    .A2(_01784_),
    .A3(_04775_),
    .B1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__o21ba_1 _12021_ (.A1(_04776_),
    .A2(_04779_),
    .B1_N(_04777_),
    .X(_05188_));
 sky130_fd_sc_hd__xnor2_2 _12022_ (.A(_05187_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__xor2_1 _12023_ (.A(_04781_),
    .B(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(_04803_),
    .B(_05190_),
    .Y(_05192_));
 sky130_fd_sc_hd__or2_1 _12025_ (.A(_04803_),
    .B(_05190_),
    .X(_05193_));
 sky130_fd_sc_hd__and2_1 _12026_ (.A(_05192_),
    .B(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__o21ai_2 _12027_ (.A1(_04783_),
    .A2(_05185_),
    .B1(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__or3_1 _12028_ (.A(_04783_),
    .B(_05185_),
    .C(_05194_),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_2 _12029_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__xor2_4 _12030_ (.A(_05184_),
    .B(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__xnor2_4 _12031_ (.A(_05183_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__a31o_2 _12032_ (.A1(_00672_),
    .A2(_03180_),
    .A3(_04800_),
    .B1(_04798_),
    .X(_05200_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_00703_),
    .B(_01251_),
    .Y(_05201_));
 sky130_fd_sc_hd__and3_2 _12034_ (.A(_01835_),
    .B(_01858_),
    .C(_05201_),
    .X(_05203_));
 sky130_fd_sc_hd__nand2_2 _12035_ (.A(_01251_),
    .B(_03180_),
    .Y(_05204_));
 sky130_fd_sc_hd__xor2_4 _12036_ (.A(_05203_),
    .B(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__xnor2_4 _12037_ (.A(_05200_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _12038_ (.A(_04357_),
    .B(_04820_),
    .Y(_05207_));
 sky130_fd_sc_hd__or2_1 _12039_ (.A(_04357_),
    .B(_04820_),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_1 _12040_ (.A(_05207_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__a21o_1 _12041_ (.A1(_04822_),
    .A2(_05209_),
    .B1(_04808_),
    .X(_05210_));
 sky130_fd_sc_hd__inv_2 _12042_ (.A(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__xnor2_4 _12043_ (.A(_05206_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_1 _12044_ (.A(_04365_),
    .B(_04830_),
    .Y(_05214_));
 sky130_fd_sc_hd__and3_1 _12045_ (.A(_04854_),
    .B(_04857_),
    .C(_04858_),
    .X(_05215_));
 sky130_fd_sc_hd__a22oi_2 _12046_ (.A1(_01250_),
    .A2(_01872_),
    .B1(_03210_),
    .B2(_01264_),
    .Y(_05216_));
 sky130_fd_sc_hd__and4_1 _12047_ (.A(_01264_),
    .B(_01250_),
    .C(_01872_),
    .D(_03210_),
    .X(_05217_));
 sky130_fd_sc_hd__a211o_1 _12048_ (.A1(_04856_),
    .A2(_04858_),
    .B1(_05216_),
    .C1(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__o211ai_1 _12049_ (.A1(_05216_),
    .A2(_05217_),
    .B1(_04856_),
    .C1(_04858_),
    .Y(_05219_));
 sky130_fd_sc_hd__and2_1 _12050_ (.A(_05218_),
    .B(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__o21a_1 _12051_ (.A1(_05215_),
    .A2(_04861_),
    .B1(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__nor3_1 _12052_ (.A(_05215_),
    .B(_04861_),
    .C(_05220_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _12053_ (.A(_05221_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_1 _12054_ (.A(_04824_),
    .B(_05223_),
    .Y(_05225_));
 sky130_fd_sc_hd__a21oi_1 _12055_ (.A1(_04827_),
    .A2(_05214_),
    .B1(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__and3_1 _12056_ (.A(_04827_),
    .B(_05214_),
    .C(_05225_),
    .X(_05227_));
 sky130_fd_sc_hd__or2_2 _12057_ (.A(_05226_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__xor2_4 _12058_ (.A(_05212_),
    .B(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__and2b_1 _12059_ (.A_N(_04831_),
    .B(_04833_),
    .X(_05230_));
 sky130_fd_sc_hd__o21ba_2 _12060_ (.A1(_04814_),
    .A2(_04834_),
    .B1_N(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__xnor2_4 _12061_ (.A(_05229_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__xnor2_4 _12062_ (.A(_05199_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _12063_ (.A(_04850_),
    .B(_04876_),
    .Y(_05234_));
 sky130_fd_sc_hd__a21bo_1 _12064_ (.A1(_04848_),
    .A2(_04877_),
    .B1_N(_05234_),
    .X(_05236_));
 sky130_fd_sc_hd__nor2_1 _12065_ (.A(_04933_),
    .B(_04935_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21bai_2 _12066_ (.A1(_04908_),
    .A2(_04936_),
    .B1_N(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__and2b_1 _12067_ (.A_N(_04872_),
    .B(_04874_),
    .X(_05239_));
 sky130_fd_sc_hd__o21ba_2 _12068_ (.A1(_04864_),
    .A2(_04875_),
    .B1_N(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_04894_),
    .B(_04903_),
    .Y(_05241_));
 sky130_fd_sc_hd__a22o_1 _12070_ (.A1(_01288_),
    .A2(_02615_),
    .B1(_02592_),
    .B2(_01309_),
    .X(_05242_));
 sky130_fd_sc_hd__inv_2 _12071_ (.A(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__and4_1 _12072_ (.A(_01309_),
    .B(_01288_),
    .C(_02615_),
    .D(_02592_),
    .X(_05244_));
 sky130_fd_sc_hd__nor2_1 _12073_ (.A(_05243_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__xnor2_2 _12074_ (.A(_04869_),
    .B(_05245_),
    .Y(_05247_));
 sky130_fd_sc_hd__or3_1 _12075_ (.A(_04867_),
    .B(_04869_),
    .C(_04870_),
    .X(_05248_));
 sky130_fd_sc_hd__a22oi_1 _12076_ (.A1(_02626_),
    .A2(_01986_),
    .B1(_03859_),
    .B2(_01365_),
    .Y(_05249_));
 sky130_fd_sc_hd__inv_2 _12077_ (.A(net216),
    .Y(_05250_));
 sky130_fd_sc_hd__or2_4 _12078_ (.A(_05250_),
    .B(_04866_),
    .X(_05251_));
 sky130_fd_sc_hd__o2111a_1 _12079_ (.A1(_00757_),
    .A2(_03859_),
    .B1(_01986_),
    .C1(_02626_),
    .D1(_01365_),
    .X(_05252_));
 sky130_fd_sc_hd__and2_1 _12080_ (.A(_05251_),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(_05249_),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__or2_1 _12082_ (.A(_05248_),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_05248_),
    .B(_05254_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05255_),
    .B(_05256_),
    .Y(_05258_));
 sky130_fd_sc_hd__xor2_2 _12085_ (.A(_05247_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__o21ai_1 _12086_ (.A1(_05241_),
    .A2(_04907_),
    .B1(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__or3_1 _12087_ (.A(_05241_),
    .B(_04907_),
    .C(_05259_),
    .X(_05261_));
 sky130_fd_sc_hd__nand2_1 _12088_ (.A(_05260_),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__xor2_2 _12089_ (.A(_05240_),
    .B(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__xor2_2 _12090_ (.A(_05238_),
    .B(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__xnor2_2 _12091_ (.A(_05236_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_04846_),
    .B(_04878_),
    .Y(_05266_));
 sky130_fd_sc_hd__a21oi_2 _12093_ (.A1(_04844_),
    .A2(_04879_),
    .B1(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__xor2_2 _12094_ (.A(_05265_),
    .B(_05267_),
    .X(_05269_));
 sky130_fd_sc_hd__xnor2_2 _12095_ (.A(_05233_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__xnor2_2 _12096_ (.A(_05181_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__xor2_2 _12097_ (.A(_05179_),
    .B(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__nand2_1 _12098_ (.A(_04965_),
    .B(_04967_),
    .Y(_05273_));
 sky130_fd_sc_hd__a21bo_1 _12099_ (.A1(_04937_),
    .A2(_04968_),
    .B1_N(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__nor2_1 _12100_ (.A(_04977_),
    .B(_05022_),
    .Y(_05275_));
 sky130_fd_sc_hd__a21o_1 _12101_ (.A1(_04975_),
    .A2(_05023_),
    .B1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__and2b_1 _12102_ (.A_N(_04916_),
    .B(_04918_),
    .X(_05277_));
 sky130_fd_sc_hd__nand2_1 _12103_ (.A(_04458_),
    .B(_04898_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(_04443_),
    .B(_04899_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _12105_ (.A(_01367_),
    .B(_02695_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_01385_),
    .B(_01367_),
    .Y(_05282_));
 sky130_fd_sc_hd__and3_1 _12107_ (.A(_02694_),
    .B(_01987_),
    .C(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__xor2_1 _12108_ (.A(_05281_),
    .B(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__a21o_1 _12109_ (.A1(_05278_),
    .A2(_05280_),
    .B1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__nand3_1 _12110_ (.A(_05278_),
    .B(_05280_),
    .C(_05284_),
    .Y(_05286_));
 sky130_fd_sc_hd__and2_1 _12111_ (.A(_05285_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _12112_ (.A1(_05277_),
    .A2(_04921_),
    .B1(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__or3_1 _12113_ (.A(_05277_),
    .B(_04921_),
    .C(_05287_),
    .X(_05289_));
 sky130_fd_sc_hd__and2_1 _12114_ (.A(_05288_),
    .B(_05289_),
    .X(_05291_));
 sky130_fd_sc_hd__or2_1 _12115_ (.A(_04901_),
    .B(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__nand2_1 _12116_ (.A(_04901_),
    .B(_05291_),
    .Y(_05293_));
 sky130_fd_sc_hd__nand2_1 _12117_ (.A(_05292_),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__o32a_1 _12118_ (.A1(_04920_),
    .A2(_04921_),
    .A3(_04932_),
    .B1(_04931_),
    .B2(_04929_),
    .X(_05295_));
 sky130_fd_sc_hd__or2b_1 _12119_ (.A(_04915_),
    .B_N(_04914_),
    .X(_05296_));
 sky130_fd_sc_hd__a22oi_1 _12120_ (.A1(_01397_),
    .A2(_02731_),
    .B1(_02019_),
    .B2(_01410_),
    .Y(_05297_));
 sky130_fd_sc_hd__and4_1 _12121_ (.A(_01410_),
    .B(_01397_),
    .C(_02731_),
    .D(_02019_),
    .X(_05298_));
 sky130_fd_sc_hd__or2_1 _12122_ (.A(_05297_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__o21ba_1 _12123_ (.A1(_04911_),
    .A2(_04913_),
    .B1_N(_04910_),
    .X(_05300_));
 sky130_fd_sc_hd__xnor2_1 _12124_ (.A(_05299_),
    .B(_05300_),
    .Y(_05302_));
 sky130_fd_sc_hd__nor2_1 _12125_ (.A(_05296_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__and2_1 _12126_ (.A(_05296_),
    .B(_05302_),
    .X(_05304_));
 sky130_fd_sc_hd__nor2_1 _12127_ (.A(_05303_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__and3_1 _12128_ (.A(_00879_),
    .B(_03967_),
    .C(_04923_),
    .X(_05306_));
 sky130_fd_sc_hd__and2b_1 _12129_ (.A_N(_04949_),
    .B(_04951_),
    .X(_05307_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(_01444_),
    .B(_03967_),
    .Y(_05308_));
 sky130_fd_sc_hd__xnor2_1 _12131_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__o21ai_1 _12132_ (.A1(_05306_),
    .A2(_04927_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__or3_1 _12133_ (.A(_05306_),
    .B(_04927_),
    .C(_05309_),
    .X(_05311_));
 sky130_fd_sc_hd__and2_1 _12134_ (.A(_05310_),
    .B(_05311_),
    .X(_05313_));
 sky130_fd_sc_hd__xor2_1 _12135_ (.A(_05305_),
    .B(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__or2b_1 _12136_ (.A(_05295_),
    .B_N(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__or2b_1 _12137_ (.A(_05314_),
    .B_N(_05295_),
    .X(_05316_));
 sky130_fd_sc_hd__nand2_1 _12138_ (.A(_05315_),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__xor2_2 _12139_ (.A(_05294_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__and2b_1 _12140_ (.A_N(_04960_),
    .B(_04946_),
    .X(_05319_));
 sky130_fd_sc_hd__a21o_1 _12141_ (.A1(_04944_),
    .A2(_04962_),
    .B1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__or2b_1 _12142_ (.A(_04996_),
    .B_N(_04999_),
    .X(_05321_));
 sky130_fd_sc_hd__o21a_1 _12143_ (.A1(_04985_),
    .A2(_05000_),
    .B1(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__and2_1 _12144_ (.A(_04952_),
    .B(_04959_),
    .X(_05324_));
 sky130_fd_sc_hd__a31o_2 _12145_ (.A1(_03999_),
    .A2(_04511_),
    .A3(_04958_),
    .B1(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__nand2_1 _12146_ (.A(_04553_),
    .B(_04980_),
    .Y(_05326_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_01443_),
    .B(_02799_),
    .Y(_05327_));
 sky130_fd_sc_hd__and3_1 _12148_ (.A(_01488_),
    .B(_02064_),
    .C(_04510_),
    .X(_05328_));
 sky130_fd_sc_hd__xnor2_1 _12149_ (.A(_05327_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__xnor2_2 _12150_ (.A(_04956_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _12151_ (.A(_00872_),
    .B(_01444_),
    .Y(_05331_));
 sky130_fd_sc_hd__and3_1 _12152_ (.A(_01434_),
    .B(_02765_),
    .C(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__xnor2_2 _12153_ (.A(_05330_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__a21oi_1 _12154_ (.A1(_05326_),
    .A2(_04984_),
    .B1(_05333_),
    .Y(_05335_));
 sky130_fd_sc_hd__and3_1 _12155_ (.A(_05326_),
    .B(_04984_),
    .C(_05333_),
    .X(_05336_));
 sky130_fd_sc_hd__nor2_1 _12156_ (.A(_05335_),
    .B(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__xnor2_1 _12157_ (.A(_05325_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__nor2_1 _12158_ (.A(_05322_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__and2_1 _12159_ (.A(_05322_),
    .B(_05338_),
    .X(_05340_));
 sky130_fd_sc_hd__nor2_1 _12160_ (.A(_05339_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__xnor2_2 _12161_ (.A(_05320_),
    .B(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__and2_1 _12162_ (.A(_04940_),
    .B(_04964_),
    .X(_05343_));
 sky130_fd_sc_hd__a21o_1 _12163_ (.A1(_04942_),
    .A2(_04963_),
    .B1(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__xor2_1 _12164_ (.A(_05342_),
    .B(_05344_),
    .X(_05346_));
 sky130_fd_sc_hd__xor2_1 _12165_ (.A(_05318_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__xnor2_1 _12166_ (.A(_05276_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__xor2_1 _12167_ (.A(_05274_),
    .B(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__a21o_1 _12168_ (.A1(_05001_),
    .A2(_05021_),
    .B1(_05019_),
    .X(_05350_));
 sky130_fd_sc_hd__nand2_1 _12169_ (.A(_05028_),
    .B(_05051_),
    .Y(_05351_));
 sky130_fd_sc_hd__a21bo_2 _12170_ (.A1(_05026_),
    .A2(_05052_),
    .B1_N(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__nor2b_1 _12171_ (.A(_04990_),
    .B_N(_04991_),
    .Y(_05353_));
 sky130_fd_sc_hd__xnor2_1 _12172_ (.A(_04539_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__a22o_1 _12173_ (.A1(_01484_),
    .A2(_02164_),
    .B1(_02132_),
    .B2(_01520_),
    .X(_05355_));
 sky130_fd_sc_hd__nand4_4 _12174_ (.A(_01520_),
    .B(_01484_),
    .C(_02164_),
    .D(_02132_),
    .Y(_05357_));
 sky130_fd_sc_hd__o21ai_1 _12175_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_04987_),
    .Y(_05358_));
 sky130_fd_sc_hd__and3_1 _12176_ (.A(_05355_),
    .B(_05357_),
    .C(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a21oi_1 _12177_ (.A1(_05355_),
    .A2(_05357_),
    .B1(_05358_),
    .Y(_05360_));
 sky130_fd_sc_hd__or2_1 _12178_ (.A(_05359_),
    .B(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__or2_1 _12179_ (.A(_04993_),
    .B(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__nand2_1 _12180_ (.A(_04993_),
    .B(_05361_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _12181_ (.A(_05362_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__or2_1 _12182_ (.A(_05354_),
    .B(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(_05354_),
    .B(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__and2_2 _12184_ (.A(_05365_),
    .B(_05366_),
    .X(_05368_));
 sky130_fd_sc_hd__nor2_1 _12185_ (.A(_05013_),
    .B(_05014_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21bo_1 _12186_ (.A1(_04612_),
    .A2(_05039_),
    .B1_N(_05037_),
    .X(_05370_));
 sky130_fd_sc_hd__and3_1 _12187_ (.A(_05007_),
    .B(_05008_),
    .C(_05010_),
    .X(_05371_));
 sky130_fd_sc_hd__a31o_1 _12188_ (.A1(_00985_),
    .A2(_03499_),
    .A3(_05011_),
    .B1(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(_00953_),
    .B(_01563_),
    .Y(_05373_));
 sky130_fd_sc_hd__and3_1 _12190_ (.A(_01524_),
    .B(_02215_),
    .C(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__nand2_1 _12191_ (.A(_01563_),
    .B(_03499_),
    .Y(_05375_));
 sky130_fd_sc_hd__xor2_1 _12192_ (.A(_05374_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__xnor2_1 _12193_ (.A(_05372_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__xor2_1 _12194_ (.A(_05370_),
    .B(_05377_),
    .X(_05379_));
 sky130_fd_sc_hd__or2_1 _12195_ (.A(_05369_),
    .B(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__nand2_1 _12196_ (.A(_05369_),
    .B(_05379_),
    .Y(_05381_));
 sky130_fd_sc_hd__and2_1 _12197_ (.A(_05380_),
    .B(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__or2b_1 _12198_ (.A(_05015_),
    .B_N(_05006_),
    .X(_05383_));
 sky130_fd_sc_hd__a21bo_1 _12199_ (.A1(_05003_),
    .A2(_05017_),
    .B1_N(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__xnor2_2 _12200_ (.A(_05382_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__xor2_2 _12201_ (.A(_05368_),
    .B(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__xnor2_2 _12202_ (.A(_05352_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__xnor2_2 _12203_ (.A(_05350_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__and3_1 _12204_ (.A(_01072_),
    .B(_03019_),
    .C(_05061_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(_01652_),
    .B(_03019_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _12206_ (.A(_01666_),
    .B(_01652_),
    .Y(_05392_));
 sky130_fd_sc_hd__and3_1 _12207_ (.A(_01667_),
    .B(_03006_),
    .C(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12208_ (.A(_05391_),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__xnor2_1 _12209_ (.A(_05390_),
    .B(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _12210_ (.A(_01629_),
    .B(_02329_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _12211_ (.A(_04659_),
    .B(_05058_),
    .Y(_05397_));
 sky130_fd_sc_hd__a21bo_1 _12212_ (.A1(_04664_),
    .A2(_05059_),
    .B1_N(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__xor2_1 _12213_ (.A(_05396_),
    .B(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__nor2_1 _12214_ (.A(_05395_),
    .B(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__and2_1 _12215_ (.A(_05395_),
    .B(_05399_),
    .X(_05402_));
 sky130_fd_sc_hd__or2_4 _12216_ (.A(_05401_),
    .B(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__and2b_1 _12217_ (.A_N(_05063_),
    .B(_05070_),
    .X(_05404_));
 sky130_fd_sc_hd__a21oi_4 _12218_ (.A1(_05054_),
    .A2(_05062_),
    .B1(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__xnor2_4 _12219_ (.A(_05403_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_05085_),
    .Y(_05407_));
 sky130_fd_sc_hd__nor2_1 _12221_ (.A(_05407_),
    .B(_05088_),
    .Y(_05408_));
 sky130_fd_sc_hd__nor2_1 _12222_ (.A(_05084_),
    .B(_05089_),
    .Y(_05409_));
 sky130_fd_sc_hd__a21bo_1 _12223_ (.A1(_05064_),
    .A2(_05065_),
    .B1_N(_05069_),
    .X(_05410_));
 sky130_fd_sc_hd__a22oi_1 _12224_ (.A1(_01603_),
    .A2(_03580_),
    .B1(_04123_),
    .B2(_01617_),
    .Y(_05412_));
 sky130_fd_sc_hd__and4_1 _12225_ (.A(_01617_),
    .B(_01603_),
    .C(_03580_),
    .D(_04123_),
    .X(_05413_));
 sky130_fd_sc_hd__or2_1 _12226_ (.A(_05412_),
    .B(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__o21ba_1 _12227_ (.A1(_04679_),
    .A2(_04681_),
    .B1_N(_05087_),
    .X(_05415_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(_01653_),
    .B(_04154_),
    .Y(_05416_));
 sky130_fd_sc_hd__mux2_2 _12229_ (.A0(_05416_),
    .A1(_04154_),
    .S(_05068_),
    .X(_05417_));
 sky130_fd_sc_hd__xor2_2 _12230_ (.A(_05415_),
    .B(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__xnor2_1 _12231_ (.A(_05414_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__or2_1 _12232_ (.A(_05410_),
    .B(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_1 _12233_ (.A(_05410_),
    .B(_05419_),
    .Y(_05421_));
 sky130_fd_sc_hd__and2_1 _12234_ (.A(_05420_),
    .B(_05421_),
    .X(_05423_));
 sky130_fd_sc_hd__o21ai_2 _12235_ (.A1(_05408_),
    .A2(_05409_),
    .B1(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__or3_1 _12236_ (.A(_05408_),
    .B(_05409_),
    .C(_05423_),
    .X(_05425_));
 sky130_fd_sc_hd__nand2_2 _12237_ (.A(_05424_),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__xor2_4 _12238_ (.A(_05406_),
    .B(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__and2b_1 _12239_ (.A_N(_05073_),
    .B(_05072_),
    .X(_05428_));
 sky130_fd_sc_hd__a21oi_2 _12240_ (.A1(_05074_),
    .A2(_05095_),
    .B1(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__xnor2_4 _12241_ (.A(_05427_),
    .B(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__o21a_2 _12242_ (.A1(_05041_),
    .A2(_05050_),
    .B1(_05047_),
    .X(_05431_));
 sky130_fd_sc_hd__and2_1 _12243_ (.A(_05078_),
    .B(_05090_),
    .X(_05432_));
 sky130_fd_sc_hd__and2_1 _12244_ (.A(_05033_),
    .B(_05035_),
    .X(_05434_));
 sky130_fd_sc_hd__a22oi_1 _12245_ (.A1(_01562_),
    .A2(_02239_),
    .B1(_02904_),
    .B2(_01584_),
    .Y(_05435_));
 sky130_fd_sc_hd__and4_1 _12246_ (.A(_01584_),
    .B(_01562_),
    .C(_02239_),
    .D(_02904_),
    .X(_05436_));
 sky130_fd_sc_hd__nor2_1 _12247_ (.A(_05435_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__o21a_1 _12248_ (.A1(_04606_),
    .A2(_05434_),
    .B1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__nor3_1 _12249_ (.A(_04606_),
    .B(_05434_),
    .C(_05437_),
    .Y(_05439_));
 sky130_fd_sc_hd__nor2_1 _12250_ (.A(_05438_),
    .B(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__nor2_1 _12251_ (.A(_05032_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__and2_1 _12252_ (.A(_05032_),
    .B(_05440_),
    .X(_05442_));
 sky130_fd_sc_hd__or2_2 _12253_ (.A(_05441_),
    .B(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__o21ai_2 _12254_ (.A1(_04639_),
    .A2(_05044_),
    .B1(_05043_),
    .Y(_05445_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(_05080_),
    .B(_05083_),
    .Y(_05446_));
 sky130_fd_sc_hd__xor2_2 _12256_ (.A(_05445_),
    .B(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__xor2_1 _12257_ (.A(_05443_),
    .B(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__o21ai_2 _12258_ (.A1(_05432_),
    .A2(_05092_),
    .B1(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__or3_1 _12259_ (.A(_05432_),
    .B(_05092_),
    .C(_05448_),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_2 _12260_ (.A(_05449_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__xor2_4 _12261_ (.A(_05431_),
    .B(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__xnor2_4 _12262_ (.A(_05430_),
    .B(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__nor2_1 _12263_ (.A(_05096_),
    .B(_05098_),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ba_2 _12264_ (.A1(_05053_),
    .A2(_05099_),
    .B1_N(_05454_),
    .X(_05456_));
 sky130_fd_sc_hd__xnor2_2 _12265_ (.A(_05453_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__xnor2_2 _12266_ (.A(_05388_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__nor2_1 _12267_ (.A(_05100_),
    .B(_05102_),
    .Y(_05459_));
 sky130_fd_sc_hd__a21oi_2 _12268_ (.A1(_05024_),
    .A2(_05103_),
    .B1(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__xor2_2 _12269_ (.A(_05458_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__xnor2_1 _12270_ (.A(_05349_),
    .B(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__nor2_1 _12271_ (.A(_05105_),
    .B(_05107_),
    .Y(_05463_));
 sky130_fd_sc_hd__a21o_1 _12272_ (.A1(_04974_),
    .A2(_05108_),
    .B1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__xnor2_1 _12273_ (.A(_05462_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__xnor2_1 _12274_ (.A(_05272_),
    .B(_05465_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _12275_ (.A(_05109_),
    .B(_05111_),
    .Y(_05468_));
 sky130_fd_sc_hd__a21oi_1 _12276_ (.A1(_04889_),
    .A2(_05112_),
    .B1(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__nor2_1 _12277_ (.A(_05467_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _12278_ (.A(_05467_),
    .B(_05469_),
    .Y(_05471_));
 sky130_fd_sc_hd__and2b_1 _12279_ (.A_N(_05470_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__xnor2_2 _12280_ (.A(_05178_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__a21oi_1 _12281_ (.A1(_04762_),
    .A2(_05118_),
    .B1(_05117_),
    .Y(_05474_));
 sky130_fd_sc_hd__xnor2_1 _12282_ (.A(_05473_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__xor2_1 _12283_ (.A(_05148_),
    .B(_05475_),
    .X(_05476_));
 sky130_fd_sc_hd__a21o_1 _12284_ (.A1(_05145_),
    .A2(_05146_),
    .B1(_05476_),
    .X(_05478_));
 sky130_fd_sc_hd__inv_2 _12285_ (.A(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__and3_1 _12286_ (.A(_05145_),
    .B(_05146_),
    .C(_05476_),
    .X(_05480_));
 sky130_fd_sc_hd__nor2_1 _12287_ (.A(_05479_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__xnor2_2 _12288_ (.A(_05144_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__xor2_2 _12289_ (.A(net262),
    .B(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__nand2_1 _12290_ (.A(_05138_),
    .B(_05142_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_1 _12291_ (.A1(_05483_),
    .A2(_05484_),
    .B1(_02185_),
    .Y(_05485_));
 sky130_fd_sc_hd__a21oi_1 _12292_ (.A1(_05483_),
    .A2(_05484_),
    .B1(_05485_),
    .Y(_00013_));
 sky130_fd_sc_hd__or2_1 _12293_ (.A(_05473_),
    .B(_05474_),
    .X(_05486_));
 sky130_fd_sc_hd__or2b_1 _12294_ (.A(_05475_),
    .B_N(_05148_),
    .X(_05488_));
 sky130_fd_sc_hd__a21o_1 _12295_ (.A1(_05150_),
    .A2(_05172_),
    .B1(_05176_),
    .X(_05489_));
 sky130_fd_sc_hd__and2b_1 _12296_ (.A_N(_05171_),
    .B(_05151_),
    .X(_05490_));
 sky130_fd_sc_hd__a21o_2 _12297_ (.A1(_05152_),
    .A2(_05170_),
    .B1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__or2b_1 _12298_ (.A(_05181_),
    .B_N(_05270_),
    .X(_05492_));
 sky130_fd_sc_hd__a21bo_1 _12299_ (.A1(_05179_),
    .A2(_05271_),
    .B1_N(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__or2b_1 _12300_ (.A(_05154_),
    .B_N(_05168_),
    .X(_05494_));
 sky130_fd_sc_hd__nand2_2 _12301_ (.A(_05166_),
    .B(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__and2b_1 _12302_ (.A_N(_05162_),
    .B(_05157_),
    .X(_05496_));
 sky130_fd_sc_hd__a31o_1 _12303_ (.A1(_01188_),
    .A2(_01754_),
    .A3(_05163_),
    .B1(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__or2b_1 _12304_ (.A(_05197_),
    .B_N(_05184_),
    .X(_05499_));
 sky130_fd_sc_hd__or2b_1 _12305_ (.A(_05198_),
    .B_N(_05183_),
    .X(_05500_));
 sky130_fd_sc_hd__nand2_1 _12306_ (.A(_02464_),
    .B(_01754_),
    .Y(_05501_));
 sky130_fd_sc_hd__and3_1 _12307_ (.A(_01157_),
    .B(_01754_),
    .C(_05159_),
    .X(_05502_));
 sky130_fd_sc_hd__a21o_1 _12308_ (.A1(_05160_),
    .A2(_05501_),
    .B1(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__a21oi_1 _12309_ (.A1(_05499_),
    .A2(_05500_),
    .B1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__and3_1 _12310_ (.A(_05499_),
    .B(_05500_),
    .C(_05503_),
    .X(_05505_));
 sky130_fd_sc_hd__nor2_1 _12311_ (.A(_05504_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__xnor2_1 _12312_ (.A(_05497_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__and2b_1 _12313_ (.A_N(_05231_),
    .B(_05229_),
    .X(_05508_));
 sky130_fd_sc_hd__a21o_1 _12314_ (.A1(_05199_),
    .A2(_05232_),
    .B1(_05508_),
    .X(_05510_));
 sky130_fd_sc_hd__or2b_1 _12315_ (.A(_05507_),
    .B_N(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__or2b_1 _12316_ (.A(_05510_),
    .B_N(_05507_),
    .X(_05512_));
 sky130_fd_sc_hd__nand2_2 _12317_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__xnor2_4 _12318_ (.A(_05495_),
    .B(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__xnor2_1 _12319_ (.A(_05493_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__xnor2_1 _12320_ (.A(_05491_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__or2b_1 _12321_ (.A(_05233_),
    .B_N(_05269_),
    .X(_05517_));
 sky130_fd_sc_hd__o21ai_2 _12322_ (.A1(_05265_),
    .A2(_05267_),
    .B1(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__and2b_1 _12323_ (.A_N(_05347_),
    .B(_05276_),
    .X(_05519_));
 sky130_fd_sc_hd__a21o_1 _12324_ (.A1(_05274_),
    .A2(_05348_),
    .B1(_05519_),
    .X(_05521_));
 sky130_fd_sc_hd__a21oi_1 _12325_ (.A1(_05206_),
    .A2(_05211_),
    .B1(_04808_),
    .Y(_05522_));
 sky130_fd_sc_hd__and2b_1 _12326_ (.A_N(_05205_),
    .B(_05200_),
    .X(_05523_));
 sky130_fd_sc_hd__nor2_1 _12327_ (.A(_05187_),
    .B(_05188_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand2_1 _12328_ (.A(_02498_),
    .B(_01784_),
    .Y(_05525_));
 sky130_fd_sc_hd__nor2_1 _12329_ (.A(_04775_),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_1 _12330_ (.A(_05524_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__inv_2 _12331_ (.A(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__xnor2_1 _12332_ (.A(_05523_),
    .B(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__o21ai_1 _12333_ (.A1(_04781_),
    .A2(_05189_),
    .B1(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__or3_1 _12334_ (.A(_04781_),
    .B(_05189_),
    .C(_05529_),
    .X(_05532_));
 sky130_fd_sc_hd__nand2_1 _12335_ (.A(_05530_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__nor2_1 _12336_ (.A(_05522_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__and2_1 _12337_ (.A(_05522_),
    .B(_05533_),
    .X(_05535_));
 sky130_fd_sc_hd__or2_1 _12338_ (.A(_05534_),
    .B(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__a21oi_2 _12339_ (.A1(_05192_),
    .A2(_05195_),
    .B1(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__and3_1 _12340_ (.A(_05192_),
    .B(_05195_),
    .C(_05536_),
    .X(_05538_));
 sky130_fd_sc_hd__nor2_2 _12341_ (.A(_05537_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__nor2_1 _12342_ (.A(_05212_),
    .B(_05228_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(_01858_),
    .B(_03180_),
    .Y(_05541_));
 sky130_fd_sc_hd__and4_2 _12344_ (.A(_01251_),
    .B(_01835_),
    .C(_01858_),
    .D(_03180_),
    .X(_05543_));
 sky130_fd_sc_hd__a21o_1 _12345_ (.A1(_04795_),
    .A2(_05541_),
    .B1(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(_05207_),
    .B(_05217_),
    .Y(_05545_));
 sky130_fd_sc_hd__xnor2_1 _12347_ (.A(_05544_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand2_1 _12348_ (.A(_01872_),
    .B(_03210_),
    .Y(_05547_));
 sky130_fd_sc_hd__a21oi_1 _12349_ (.A1(_04869_),
    .A2(_05242_),
    .B1(_05244_),
    .Y(_05548_));
 sky130_fd_sc_hd__xnor2_1 _12350_ (.A(_05547_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__and2_1 _12351_ (.A(_05218_),
    .B(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__nor2_1 _12352_ (.A(_05218_),
    .B(_05549_),
    .Y(_05551_));
 sky130_fd_sc_hd__nor2_1 _12353_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__a21o_1 _12354_ (.A1(_04824_),
    .A2(_05223_),
    .B1(_05221_),
    .X(_05554_));
 sky130_fd_sc_hd__and2_1 _12355_ (.A(_05552_),
    .B(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__nor2_1 _12356_ (.A(_05552_),
    .B(_05554_),
    .Y(_05556_));
 sky130_fd_sc_hd__nor2_1 _12357_ (.A(_05555_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__xnor2_1 _12358_ (.A(_05546_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__o21a_1 _12359_ (.A1(_05226_),
    .A2(_05540_),
    .B1(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__nor3_1 _12360_ (.A(_05226_),
    .B(_05540_),
    .C(_05558_),
    .Y(_05560_));
 sky130_fd_sc_hd__nor2_2 _12361_ (.A(_05559_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__xnor2_4 _12362_ (.A(_05539_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__o21ai_2 _12363_ (.A1(_05240_),
    .A2(_05262_),
    .B1(_05260_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21a_1 _12364_ (.A1(_05294_),
    .A2(_05317_),
    .B1(_05315_),
    .X(_05565_));
 sky130_fd_sc_hd__o21a_2 _12365_ (.A1(_05247_),
    .A2(_05258_),
    .B1(_05255_),
    .X(_05566_));
 sky130_fd_sc_hd__nand2_1 _12366_ (.A(_05288_),
    .B(_05293_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand2_2 _12367_ (.A(_02615_),
    .B(_02592_),
    .Y(_05568_));
 sky130_fd_sc_hd__xnor2_4 _12368_ (.A(_05251_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _12369_ (.A(_01986_),
    .B(_03859_),
    .Y(_05570_));
 sky130_fd_sc_hd__mux2_4 _12370_ (.A0(_05570_),
    .A1(_03859_),
    .S(_05253_),
    .X(_05571_));
 sky130_fd_sc_hd__xnor2_4 _12371_ (.A(_05569_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__xor2_2 _12372_ (.A(_05567_),
    .B(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__xor2_2 _12373_ (.A(_05566_),
    .B(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__xnor2_2 _12374_ (.A(_05565_),
    .B(_05574_),
    .Y(_05576_));
 sky130_fd_sc_hd__xnor2_2 _12375_ (.A(_05563_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__and2_1 _12376_ (.A(_05238_),
    .B(_05263_),
    .X(_05578_));
 sky130_fd_sc_hd__a21oi_2 _12377_ (.A1(_05236_),
    .A2(_05264_),
    .B1(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__xor2_2 _12378_ (.A(_05577_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__xnor2_2 _12379_ (.A(_05562_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_1 _12380_ (.A(_05521_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__xnor2_1 _12381_ (.A(_05518_),
    .B(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__inv_2 _12382_ (.A(_05346_),
    .Y(_05584_));
 sky130_fd_sc_hd__or2b_1 _12383_ (.A(_05342_),
    .B_N(_05344_),
    .X(_05585_));
 sky130_fd_sc_hd__a21bo_1 _12384_ (.A1(_05318_),
    .A2(_05584_),
    .B1_N(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__and2b_1 _12385_ (.A_N(_05386_),
    .B(_05352_),
    .X(_05588_));
 sky130_fd_sc_hd__a21o_1 _12386_ (.A1(_05350_),
    .A2(_05387_),
    .B1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__inv_2 _12387_ (.A(_02695_),
    .Y(_05590_));
 sky130_fd_sc_hd__a31o_1 _12388_ (.A1(_01385_),
    .A2(_02694_),
    .A3(_01367_),
    .B1(_02695_),
    .X(_05591_));
 sky130_fd_sc_hd__o211a_1 _12389_ (.A1(_05590_),
    .A2(_04897_),
    .B1(_05591_),
    .C1(_01987_),
    .X(_05592_));
 sky130_fd_sc_hd__xnor2_1 _12390_ (.A(_05303_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__and2_1 _12391_ (.A(_05285_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__nor2_1 _12392_ (.A(_05285_),
    .B(_05593_),
    .Y(_05595_));
 sky130_fd_sc_hd__or2_1 _12393_ (.A(_05594_),
    .B(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__nor2_1 _12394_ (.A(_05299_),
    .B(_05300_),
    .Y(_05598_));
 sky130_fd_sc_hd__nand2_1 _12395_ (.A(_01410_),
    .B(_01397_),
    .Y(_05599_));
 sky130_fd_sc_hd__and3_1 _12396_ (.A(_02731_),
    .B(_02019_),
    .C(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__nand2_2 _12397_ (.A(_05598_),
    .B(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__or2_1 _12398_ (.A(_05598_),
    .B(_05600_),
    .X(_05602_));
 sky130_fd_sc_hd__nand2_1 _12399_ (.A(_05601_),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__or3b_1 _12400_ (.A(_04949_),
    .B(_05308_),
    .C_N(_04951_),
    .X(_05604_));
 sky130_fd_sc_hd__nand2_1 _12401_ (.A(_02765_),
    .B(_03967_),
    .Y(_05605_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(_05605_),
    .A1(_03967_),
    .S(_04948_),
    .X(_05606_));
 sky130_fd_sc_hd__or2_1 _12403_ (.A(_05604_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__nand2_1 _12404_ (.A(_05604_),
    .B(_05606_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _12405_ (.A(_05607_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__or2_1 _12406_ (.A(_05603_),
    .B(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__nand2_1 _12407_ (.A(_05603_),
    .B(_05610_),
    .Y(_05612_));
 sky130_fd_sc_hd__and2_1 _12408_ (.A(_05611_),
    .B(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__a21bo_1 _12409_ (.A1(_05305_),
    .A2(_05311_),
    .B1_N(_05310_),
    .X(_05614_));
 sky130_fd_sc_hd__xnor2_1 _12410_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__nor2_1 _12411_ (.A(_05596_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(_05596_),
    .B(_05615_),
    .Y(_05617_));
 sky130_fd_sc_hd__or2b_2 _12413_ (.A(_05616_),
    .B_N(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__a21oi_2 _12414_ (.A1(_05320_),
    .A2(_05341_),
    .B1(_05339_),
    .Y(_05620_));
 sky130_fd_sc_hd__a21oi_2 _12415_ (.A1(_05325_),
    .A2(_05337_),
    .B1(_05335_),
    .Y(_05621_));
 sky130_fd_sc_hd__or4_1 _12416_ (.A(_04509_),
    .B(_04510_),
    .C(_04954_),
    .D(_05327_),
    .X(_05622_));
 sky130_fd_sc_hd__a21bo_1 _12417_ (.A1(_05330_),
    .A2(_05332_),
    .B1_N(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__inv_2 _12418_ (.A(_01487_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_1 _12419_ (.A1(_05624_),
    .A2(_02799_),
    .B1(_04953_),
    .Y(_05625_));
 sky130_fd_sc_hd__o211a_1 _12420_ (.A1(_02799_),
    .A2(_04953_),
    .B1(_05625_),
    .C1(_02064_),
    .X(_05626_));
 sky130_fd_sc_hd__and3_1 _12421_ (.A(_04539_),
    .B(_05353_),
    .C(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__a21oi_1 _12422_ (.A1(_04539_),
    .A2(_05353_),
    .B1(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__nor2_1 _12423_ (.A(_05627_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__xnor2_1 _12424_ (.A(_05623_),
    .B(_05629_),
    .Y(_05631_));
 sky130_fd_sc_hd__a21oi_1 _12425_ (.A1(_05362_),
    .A2(_05365_),
    .B1(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__and3_1 _12426_ (.A(_05362_),
    .B(_05365_),
    .C(_05631_),
    .X(_05633_));
 sky130_fd_sc_hd__nor2_1 _12427_ (.A(_05632_),
    .B(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__xnor2_2 _12428_ (.A(_05621_),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__and2b_1 _12429_ (.A_N(_05620_),
    .B(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__and2b_1 _12430_ (.A_N(_05635_),
    .B(_05620_),
    .X(_05637_));
 sky130_fd_sc_hd__nor2_1 _12431_ (.A(_05636_),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__xnor2_1 _12432_ (.A(_05618_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__xnor2_1 _12433_ (.A(_05589_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__xnor2_1 _12434_ (.A(_05587_),
    .B(_05640_),
    .Y(_05642_));
 sky130_fd_sc_hd__and2_1 _12435_ (.A(_05390_),
    .B(_05394_),
    .X(_05643_));
 sky130_fd_sc_hd__inv_2 _12436_ (.A(_03019_),
    .Y(_05644_));
 sky130_fd_sc_hd__a31o_1 _12437_ (.A1(_01666_),
    .A2(_01667_),
    .A3(_01652_),
    .B1(_03019_),
    .X(_05645_));
 sky130_fd_sc_hd__o211a_1 _12438_ (.A1(_05644_),
    .A2(_05057_),
    .B1(_05645_),
    .C1(_03006_),
    .X(_05646_));
 sky130_fd_sc_hd__o21a_1 _12439_ (.A1(_05643_),
    .A2(_05401_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nor3_1 _12440_ (.A(_05643_),
    .B(_05401_),
    .C(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__nor2_2 _12441_ (.A(_05647_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__o32ai_4 _12442_ (.A1(_05086_),
    .A2(_05087_),
    .A3(_05417_),
    .B1(_05418_),
    .B2(_05414_),
    .Y(_05650_));
 sky130_fd_sc_hd__and3_1 _12443_ (.A(_01629_),
    .B(_02329_),
    .C(_05398_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2_1 _12444_ (.A(_03580_),
    .B(_04123_),
    .Y(_05653_));
 sky130_fd_sc_hd__and3b_1 _12445_ (.A_N(_05068_),
    .B(_04154_),
    .C(_02329_),
    .X(_05654_));
 sky130_fd_sc_hd__xnor2_1 _12446_ (.A(_05653_),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_1 _12447_ (.A(_05651_),
    .B(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__nor2_1 _12448_ (.A(_05651_),
    .B(_05655_),
    .Y(_05657_));
 sky130_fd_sc_hd__or2_1 _12449_ (.A(_05656_),
    .B(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__xnor2_2 _12450_ (.A(_05650_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__xor2_4 _12451_ (.A(_05649_),
    .B(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__or2_1 _12452_ (.A(_05406_),
    .B(_05426_),
    .X(_05661_));
 sky130_fd_sc_hd__o21ai_4 _12453_ (.A1(_05403_),
    .A2(_05405_),
    .B1(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_4 _12454_ (.A(_05660_),
    .B(_05662_),
    .Y(_05664_));
 sky130_fd_sc_hd__or2b_1 _12455_ (.A(_05445_),
    .B_N(_05446_),
    .X(_05665_));
 sky130_fd_sc_hd__o21ai_4 _12456_ (.A1(_05443_),
    .A2(_05447_),
    .B1(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _12457_ (.A(_01584_),
    .B(_01562_),
    .Y(_05667_));
 sky130_fd_sc_hd__and4_1 _12458_ (.A(_02239_),
    .B(_02904_),
    .C(_05667_),
    .D(_05413_),
    .X(_05668_));
 sky130_fd_sc_hd__a31o_1 _12459_ (.A1(_02239_),
    .A2(_02904_),
    .A3(_05667_),
    .B1(_05413_),
    .X(_05669_));
 sky130_fd_sc_hd__or2b_1 _12460_ (.A(_05668_),
    .B_N(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__a21oi_1 _12461_ (.A1(_05420_),
    .A2(_05424_),
    .B1(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__and3_1 _12462_ (.A(_05420_),
    .B(_05424_),
    .C(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nor2_2 _12463_ (.A(_05671_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_4 _12464_ (.A(_05666_),
    .B(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__xnor2_4 _12465_ (.A(_05664_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__and2b_1 _12466_ (.A_N(_05429_),
    .B(_05427_),
    .X(_05677_));
 sky130_fd_sc_hd__a21oi_4 _12467_ (.A1(_05430_),
    .A2(_05452_),
    .B1(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__xnor2_2 _12468_ (.A(_05676_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__inv_2 _12469_ (.A(_05385_),
    .Y(_05680_));
 sky130_fd_sc_hd__a32o_1 _12470_ (.A1(_05380_),
    .A2(_05381_),
    .A3(_05384_),
    .B1(_05680_),
    .B2(_05368_),
    .X(_05681_));
 sky130_fd_sc_hd__o21ai_4 _12471_ (.A1(_05431_),
    .A2(_05451_),
    .B1(_05449_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_1 _12472_ (.A(_01520_),
    .B(_01484_),
    .Y(_05683_));
 sky130_fd_sc_hd__and3_1 _12473_ (.A(_02164_),
    .B(_02132_),
    .C(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__nand2_1 _12474_ (.A(_05359_),
    .B(_05684_),
    .Y(_05686_));
 sky130_fd_sc_hd__or2_1 _12475_ (.A(_05359_),
    .B(_05684_),
    .X(_05687_));
 sky130_fd_sc_hd__nand2_2 _12476_ (.A(_05686_),
    .B(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_05370_),
    .B(_05377_),
    .Y(_05689_));
 sky130_fd_sc_hd__and2b_1 _12478_ (.A_N(_05376_),
    .B(_05372_),
    .X(_05690_));
 sky130_fd_sc_hd__nand2_1 _12479_ (.A(_02215_),
    .B(_03499_),
    .Y(_05691_));
 sky130_fd_sc_hd__and4_1 _12480_ (.A(_01563_),
    .B(_01524_),
    .C(_02215_),
    .D(_03499_),
    .X(_05692_));
 sky130_fd_sc_hd__a21oi_1 _12481_ (.A1(_05008_),
    .A2(_05691_),
    .B1(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_2 _12482_ (.A1(_05438_),
    .A2(_05442_),
    .B1(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__or3_1 _12483_ (.A(_05438_),
    .B(_05442_),
    .C(_05693_),
    .X(_05695_));
 sky130_fd_sc_hd__and2_1 _12484_ (.A(_05694_),
    .B(_05695_),
    .X(_05697_));
 sky130_fd_sc_hd__xnor2_1 _12485_ (.A(_05690_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__a21o_1 _12486_ (.A1(_05689_),
    .A2(_05381_),
    .B1(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__nand3_1 _12487_ (.A(_05689_),
    .B(_05381_),
    .C(_05698_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(_05699_),
    .B(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__xor2_2 _12489_ (.A(_05688_),
    .B(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__xor2_2 _12490_ (.A(_05682_),
    .B(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__xor2_2 _12491_ (.A(_05681_),
    .B(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__xnor2_2 _12492_ (.A(_05679_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__or2_1 _12493_ (.A(_05453_),
    .B(_05456_),
    .X(_05706_));
 sky130_fd_sc_hd__o21a_1 _12494_ (.A1(_05388_),
    .A2(_05457_),
    .B1(_05706_),
    .X(_05708_));
 sky130_fd_sc_hd__xnor2_2 _12495_ (.A(_05705_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__xnor2_1 _12496_ (.A(_05642_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__nor2_1 _12497_ (.A(_05458_),
    .B(_05460_),
    .Y(_05711_));
 sky130_fd_sc_hd__a21oi_1 _12498_ (.A1(_05349_),
    .A2(_05461_),
    .B1(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__xor2_1 _12499_ (.A(_05710_),
    .B(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__xnor2_1 _12500_ (.A(_05583_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__or2b_1 _12501_ (.A(_05462_),
    .B_N(_05464_),
    .X(_05715_));
 sky130_fd_sc_hd__a21boi_1 _12502_ (.A1(_05272_),
    .A2(_05465_),
    .B1_N(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__nor2_1 _12503_ (.A(_05714_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_1 _12504_ (.A(_05714_),
    .B(_05716_),
    .Y(_05719_));
 sky130_fd_sc_hd__and2b_1 _12505_ (.A_N(_05717_),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__xnor2_1 _12506_ (.A(_05516_),
    .B(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__a21oi_1 _12507_ (.A1(_05178_),
    .A2(_05471_),
    .B1(_05470_),
    .Y(_05722_));
 sky130_fd_sc_hd__nor2_1 _12508_ (.A(_05721_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__and2_1 _12509_ (.A(_05721_),
    .B(_05722_),
    .X(_05724_));
 sky130_fd_sc_hd__nor2_1 _12510_ (.A(_05723_),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__xnor2_2 _12511_ (.A(_05489_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__a21oi_2 _12512_ (.A1(_05486_),
    .A2(_05488_),
    .B1(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__and3_1 _12513_ (.A(_05486_),
    .B(_05488_),
    .C(_05726_),
    .X(_05728_));
 sky130_fd_sc_hd__nor2_2 _12514_ (.A(_05727_),
    .B(_05728_),
    .Y(_05730_));
 sky130_fd_sc_hd__a21o_1 _12515_ (.A1(_05128_),
    .A2(_05478_),
    .B1(_05480_),
    .X(_05731_));
 sky130_fd_sc_hd__inv_2 _12516_ (.A(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__a31o_4 _12517_ (.A1(_05130_),
    .A2(_05135_),
    .A3(_05481_),
    .B1(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__xor2_2 _12518_ (.A(_05730_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__xor2_1 _12519_ (.A(net263),
    .B(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__a21oi_1 _12520_ (.A1(_04243_),
    .A2(_04726_),
    .B1(_04722_),
    .Y(_05736_));
 sky130_fd_sc_hd__a41o_1 _12521_ (.A1(_03691_),
    .A2(_03692_),
    .A3(_04245_),
    .A4(_04723_),
    .B1(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__and3_1 _12522_ (.A(_05138_),
    .B(_05139_),
    .C(_05483_),
    .X(_05738_));
 sky130_fd_sc_hd__nand2_1 _12523_ (.A(net262),
    .B(_05482_),
    .Y(_05739_));
 sky130_fd_sc_hd__nor2_1 _12524_ (.A(net262),
    .B(_05482_),
    .Y(_05741_));
 sky130_fd_sc_hd__a21oi_1 _12525_ (.A1(_05138_),
    .A2(_05739_),
    .B1(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__a21o_1 _12526_ (.A1(_05737_),
    .A2(_05738_),
    .B1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(_05735_),
    .B(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_05735_),
    .B(_05743_),
    .Y(_05745_));
 sky130_fd_sc_hd__and3_1 _12529_ (.A(_02174_),
    .B(_05744_),
    .C(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__clkbuf_1 _12530_ (.A(_05746_),
    .X(_00014_));
 sky130_fd_sc_hd__a21oi_4 _12531_ (.A1(_05730_),
    .A2(_05733_),
    .B1(_05727_),
    .Y(_05747_));
 sky130_fd_sc_hd__or2b_1 _12532_ (.A(_05515_),
    .B_N(_05491_),
    .X(_05748_));
 sky130_fd_sc_hd__a21bo_2 _12533_ (.A1(_05493_),
    .A2(_05514_),
    .B1_N(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__or2b_1 _12534_ (.A(_05513_),
    .B_N(_05495_),
    .X(_05751_));
 sky130_fd_sc_hd__nand2_2 _12535_ (.A(_05511_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__or2b_1 _12536_ (.A(_05582_),
    .B_N(_05518_),
    .X(_05753_));
 sky130_fd_sc_hd__a21bo_1 _12537_ (.A1(_05521_),
    .A2(_05581_),
    .B1_N(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__a21o_1 _12538_ (.A1(_05497_),
    .A2(_05506_),
    .B1(_05504_),
    .X(_05755_));
 sky130_fd_sc_hd__a21o_1 _12539_ (.A1(_05539_),
    .A2(_05561_),
    .B1(_05559_),
    .X(_05756_));
 sky130_fd_sc_hd__o21a_2 _12540_ (.A1(_05534_),
    .A2(_05537_),
    .B1(_05502_),
    .X(_05757_));
 sky130_fd_sc_hd__nor3_1 _12541_ (.A(_05502_),
    .B(_05534_),
    .C(_05537_),
    .Y(_05758_));
 sky130_fd_sc_hd__nor2_1 _12542_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__xor2_1 _12543_ (.A(_05756_),
    .B(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__and2_1 _12544_ (.A(_05755_),
    .B(_05760_),
    .X(_05762_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(_05755_),
    .B(_05760_),
    .Y(_05763_));
 sky130_fd_sc_hd__nor2_2 _12546_ (.A(_05762_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__xnor2_1 _12547_ (.A(_05754_),
    .B(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__xnor2_1 _12548_ (.A(_05752_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__or2b_1 _12549_ (.A(_05562_),
    .B_N(_05580_),
    .X(_05767_));
 sky130_fd_sc_hd__o21ai_2 _12550_ (.A1(_05577_),
    .A2(_05579_),
    .B1(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__or2b_1 _12551_ (.A(_05640_),
    .B_N(_05587_),
    .X(_05769_));
 sky130_fd_sc_hd__a21bo_1 _12552_ (.A1(_05589_),
    .A2(_05639_),
    .B1_N(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a21bo_1 _12553_ (.A1(_05523_),
    .A2(_05528_),
    .B1_N(_05532_),
    .X(_05771_));
 sky130_fd_sc_hd__o21ai_2 _12554_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05207_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21ba_1 _12555_ (.A1(_04775_),
    .A2(_05524_),
    .B1_N(_05525_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_2 _12556_ (.A(_05543_),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(_05543_),
    .B(_05774_),
    .X(_05776_));
 sky130_fd_sc_hd__and2_1 _12558_ (.A(_05775_),
    .B(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__nand2_1 _12559_ (.A(_05773_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__or2_1 _12560_ (.A(_05773_),
    .B(_05777_),
    .X(_05779_));
 sky130_fd_sc_hd__and2_1 _12561_ (.A(_05778_),
    .B(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__xor2_1 _12562_ (.A(_05771_),
    .B(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(_05552_),
    .B(_05554_),
    .Y(_05782_));
 sky130_fd_sc_hd__o21a_1 _12564_ (.A1(_05546_),
    .A2(_05556_),
    .B1(_05782_),
    .X(_05784_));
 sky130_fd_sc_hd__a41o_1 _12565_ (.A1(_01872_),
    .A2(_03210_),
    .A3(_04869_),
    .A4(_05245_),
    .B1(_05551_),
    .X(_05785_));
 sky130_fd_sc_hd__nand3_1 _12566_ (.A(_01872_),
    .B(_03210_),
    .C(_05244_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_1 _12567_ (.A1(_05251_),
    .A2(_05568_),
    .B1(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21a_1 _12568_ (.A1(_05251_),
    .A2(_05786_),
    .B1(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__xor2_1 _12569_ (.A(_05785_),
    .B(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__and2b_2 _12570_ (.A_N(_05784_),
    .B(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__and2b_1 _12571_ (.A_N(_05789_),
    .B(_05784_),
    .X(_05791_));
 sky130_fd_sc_hd__nor2_2 _12572_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__and2_1 _12573_ (.A(_05781_),
    .B(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__nor2_1 _12574_ (.A(_05781_),
    .B(_05792_),
    .Y(_05795_));
 sky130_fd_sc_hd__nor2_2 _12575_ (.A(_05793_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21o_1 _12576_ (.A1(_05288_),
    .A2(_05293_),
    .B1(_05572_),
    .X(_05797_));
 sky130_fd_sc_hd__o21ai_2 _12577_ (.A1(_05566_),
    .A2(_05573_),
    .B1(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__and2_1 _12578_ (.A(_05613_),
    .B(_05614_),
    .X(_05799_));
 sky130_fd_sc_hd__a21oi_1 _12579_ (.A1(_05303_),
    .A2(_05592_),
    .B1(_05595_),
    .Y(_05800_));
 sky130_fd_sc_hd__o2bb2ai_4 _12580_ (.A1_N(_03859_),
    .A2_N(_05253_),
    .B1(_05569_),
    .B2(_05571_),
    .Y(_05801_));
 sky130_fd_sc_hd__xnor2_1 _12581_ (.A(_05800_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_1 _12582_ (.A1(_05799_),
    .A2(_05616_),
    .B1(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__or3_1 _12583_ (.A(_05799_),
    .B(_05616_),
    .C(_05802_),
    .X(_05804_));
 sky130_fd_sc_hd__and2_1 _12584_ (.A(_05803_),
    .B(_05804_),
    .X(_05806_));
 sky130_fd_sc_hd__xnor2_1 _12585_ (.A(_05798_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__and2b_1 _12586_ (.A_N(_05565_),
    .B(_05574_),
    .X(_05808_));
 sky130_fd_sc_hd__a21oi_1 _12587_ (.A1(_05563_),
    .A2(_05576_),
    .B1(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nor2_1 _12588_ (.A(_05807_),
    .B(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__and2_1 _12589_ (.A(_05807_),
    .B(_05809_),
    .X(_05811_));
 sky130_fd_sc_hd__nor2_1 _12590_ (.A(_05810_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__xnor2_1 _12591_ (.A(_05796_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__xnor2_1 _12592_ (.A(_05770_),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__xnor2_1 _12593_ (.A(_05768_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__nor2_1 _12594_ (.A(_05676_),
    .B(_05678_),
    .Y(_05817_));
 sky130_fd_sc_hd__and2b_1 _12595_ (.A_N(_05679_),
    .B(_05704_),
    .X(_05818_));
 sky130_fd_sc_hd__and4_1 _12596_ (.A(_01667_),
    .B(_01652_),
    .C(_03019_),
    .D(_03006_),
    .X(_05819_));
 sky130_fd_sc_hd__a32o_1 _12597_ (.A1(_03580_),
    .A2(_04123_),
    .A3(_05654_),
    .B1(_05068_),
    .B2(_04154_),
    .X(_05820_));
 sky130_fd_sc_hd__nand2_1 _12598_ (.A(_05819_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__or2_1 _12599_ (.A(_05819_),
    .B(_05820_),
    .X(_05822_));
 sky130_fd_sc_hd__and2_1 _12600_ (.A(_05821_),
    .B(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__a21o_1 _12601_ (.A1(_05649_),
    .A2(_05659_),
    .B1(_05647_),
    .X(_05824_));
 sky130_fd_sc_hd__xor2_1 _12602_ (.A(_05823_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__and2b_1 _12603_ (.A_N(_05658_),
    .B(_05650_),
    .X(_05826_));
 sky130_fd_sc_hd__o21a_1 _12604_ (.A1(_05656_),
    .A2(_05826_),
    .B1(_05668_),
    .X(_05828_));
 sky130_fd_sc_hd__nor3_1 _12605_ (.A(_05656_),
    .B(_05826_),
    .C(_05668_),
    .Y(_05829_));
 sky130_fd_sc_hd__nor2_1 _12606_ (.A(_05828_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_1 _12607_ (.A(_05825_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__or2_1 _12608_ (.A(_05825_),
    .B(_05830_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _12609_ (.A(_05831_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _12610_ (.A(_05660_),
    .B(_05662_),
    .Y(_05834_));
 sky130_fd_sc_hd__o21a_2 _12611_ (.A1(_05664_),
    .A2(_05675_),
    .B1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__xnor2_1 _12612_ (.A(_05833_),
    .B(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__o21a_1 _12613_ (.A1(_05688_),
    .A2(_05701_),
    .B1(_05699_),
    .X(_05837_));
 sky130_fd_sc_hd__a21o_2 _12614_ (.A1(_05666_),
    .A2(_05673_),
    .B1(_05671_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _12615_ (.A(_05690_),
    .B(_05697_),
    .Y(_05840_));
 sky130_fd_sc_hd__xnor2_1 _12616_ (.A(_05436_),
    .B(_05692_),
    .Y(_05841_));
 sky130_fd_sc_hd__a21o_1 _12617_ (.A1(_05694_),
    .A2(_05840_),
    .B1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__nand3_1 _12618_ (.A(_05694_),
    .B(_05840_),
    .C(_05841_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_1 _12619_ (.A(_05842_),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__xnor2_2 _12620_ (.A(_05357_),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__xnor2_2 _12621_ (.A(_05839_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__xnor2_2 _12622_ (.A(_05837_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_1 _12623_ (.A(_05836_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21a_1 _12624_ (.A1(_05817_),
    .A2(_05818_),
    .B1(_05848_),
    .X(_05850_));
 sky130_fd_sc_hd__nor3_1 _12625_ (.A(_05817_),
    .B(_05818_),
    .C(_05848_),
    .Y(_05851_));
 sky130_fd_sc_hd__nor2_1 _12626_ (.A(_05850_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ba_1 _12627_ (.A1(_05618_),
    .A2(_05637_),
    .B1_N(_05636_),
    .X(_05853_));
 sky130_fd_sc_hd__and2_1 _12628_ (.A(_05682_),
    .B(_05702_),
    .X(_05854_));
 sky130_fd_sc_hd__and2_1 _12629_ (.A(_05681_),
    .B(_05703_),
    .X(_05855_));
 sky130_fd_sc_hd__and4_1 _12630_ (.A(_02694_),
    .B(_01367_),
    .C(_02695_),
    .D(_01987_),
    .X(_05856_));
 sky130_fd_sc_hd__xor2_2 _12631_ (.A(_05601_),
    .B(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__and3_2 _12632_ (.A(_03967_),
    .B(_04948_),
    .C(_05298_),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_1 _12633_ (.A1(_03967_),
    .A2(_04948_),
    .B1(_05298_),
    .Y(_05859_));
 sky130_fd_sc_hd__or2_1 _12634_ (.A(_05858_),
    .B(_05859_),
    .X(_05861_));
 sky130_fd_sc_hd__a21o_1 _12635_ (.A1(_05607_),
    .A2(_05611_),
    .B1(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__nand3_1 _12636_ (.A(_05607_),
    .B(_05611_),
    .C(_05861_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _12637_ (.A(_05862_),
    .B(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__xnor2_2 _12638_ (.A(_05857_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_1 _12639_ (.A1(_05623_),
    .A2(_05629_),
    .B1(_05627_),
    .X(_05866_));
 sky130_fd_sc_hd__and4_2 _12640_ (.A(_01488_),
    .B(_01443_),
    .C(_02799_),
    .D(_02064_),
    .X(_05867_));
 sky130_fd_sc_hd__xnor2_1 _12641_ (.A(_05686_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__and2_1 _12642_ (.A(_05866_),
    .B(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__or2_1 _12643_ (.A(_05866_),
    .B(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__or2b_1 _12644_ (.A(_05869_),
    .B_N(_05870_),
    .X(_05872_));
 sky130_fd_sc_hd__o21ba_1 _12645_ (.A1(_05621_),
    .A2(_05633_),
    .B1_N(_05632_),
    .X(_05873_));
 sky130_fd_sc_hd__nor2_1 _12646_ (.A(_05872_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__and2_1 _12647_ (.A(_05872_),
    .B(_05873_),
    .X(_05875_));
 sky130_fd_sc_hd__or2_1 _12648_ (.A(_05874_),
    .B(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__xor2_1 _12649_ (.A(_05865_),
    .B(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__o21a_1 _12650_ (.A1(_05854_),
    .A2(_05855_),
    .B1(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__nor3_1 _12651_ (.A(_05854_),
    .B(_05855_),
    .C(_05877_),
    .Y(_05879_));
 sky130_fd_sc_hd__nor2_1 _12652_ (.A(_05878_),
    .B(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__xnor2_2 _12653_ (.A(_05853_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__xnor2_1 _12654_ (.A(_05852_),
    .B(_05881_),
    .Y(_05883_));
 sky130_fd_sc_hd__and2b_1 _12655_ (.A_N(_05708_),
    .B(_05705_),
    .X(_05884_));
 sky130_fd_sc_hd__a21o_1 _12656_ (.A1(_05642_),
    .A2(_05709_),
    .B1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__xor2_1 _12657_ (.A(_05883_),
    .B(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__xnor2_1 _12658_ (.A(_05815_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nor2_1 _12659_ (.A(_05710_),
    .B(_05712_),
    .Y(_05888_));
 sky130_fd_sc_hd__a21oi_1 _12660_ (.A1(_05583_),
    .A2(_05713_),
    .B1(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__xor2_1 _12661_ (.A(_05887_),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__xnor2_1 _12662_ (.A(_05766_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__a21oi_1 _12663_ (.A1(_05516_),
    .A2(_05719_),
    .B1(_05717_),
    .Y(_05892_));
 sky130_fd_sc_hd__nor2_1 _12664_ (.A(_05891_),
    .B(_05892_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_1 _12665_ (.A(_05891_),
    .B(_05892_),
    .Y(_05895_));
 sky130_fd_sc_hd__and2b_1 _12666_ (.A_N(_05894_),
    .B(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__xnor2_4 _12667_ (.A(_05749_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__a21o_1 _12668_ (.A1(_05489_),
    .A2(_05725_),
    .B1(_05723_),
    .X(_05898_));
 sky130_fd_sc_hd__xnor2_2 _12669_ (.A(_05897_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__xnor2_2 _12670_ (.A(_05747_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__xor2_2 _12671_ (.A(net264),
    .B(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__a21bo_1 _12672_ (.A1(net263),
    .A2(_05734_),
    .B1_N(_05745_),
    .X(_05902_));
 sky130_fd_sc_hd__o21ai_1 _12673_ (.A1(_05901_),
    .A2(_05902_),
    .B1(_02185_),
    .Y(_05903_));
 sky130_fd_sc_hd__a21oi_1 _12674_ (.A1(_05901_),
    .A2(_05902_),
    .B1(_05903_),
    .Y(_00015_));
 sky130_fd_sc_hd__o21a_1 _12675_ (.A1(_05357_),
    .A2(_05844_),
    .B1(_05842_),
    .X(_05905_));
 sky130_fd_sc_hd__a21oi_2 _12676_ (.A1(_05436_),
    .A2(_05692_),
    .B1(_05828_),
    .Y(_05906_));
 sky130_fd_sc_hd__xnor2_2 _12677_ (.A(_05905_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__xor2_1 _12678_ (.A(_05821_),
    .B(_05831_),
    .X(_05908_));
 sky130_fd_sc_hd__a21oi_2 _12679_ (.A1(_05823_),
    .A2(_05824_),
    .B1(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__xor2_2 _12680_ (.A(_05907_),
    .B(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__nand2_1 _12681_ (.A(_05833_),
    .B(_05835_),
    .Y(_05911_));
 sky130_fd_sc_hd__nor2_1 _12682_ (.A(_05833_),
    .B(_05835_),
    .Y(_05912_));
 sky130_fd_sc_hd__a21oi_2 _12683_ (.A1(_05911_),
    .A2(_05847_),
    .B1(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_1 _12684_ (.A(_05910_),
    .B(_05913_),
    .Y(_05915_));
 sky130_fd_sc_hd__o21ba_1 _12685_ (.A1(_05865_),
    .A2(_05876_),
    .B1_N(_05874_),
    .X(_05916_));
 sky130_fd_sc_hd__and2b_1 _12686_ (.A_N(_05845_),
    .B(_05839_),
    .X(_05917_));
 sky130_fd_sc_hd__and2b_1 _12687_ (.A_N(_05837_),
    .B(_05846_),
    .X(_05918_));
 sky130_fd_sc_hd__and3_1 _12688_ (.A(_05359_),
    .B(_05684_),
    .C(_05867_),
    .X(_05919_));
 sky130_fd_sc_hd__o21ai_4 _12689_ (.A1(_05919_),
    .A2(_05869_),
    .B1(_05858_),
    .Y(_05920_));
 sky130_fd_sc_hd__or3_1 _12690_ (.A(_05858_),
    .B(_05919_),
    .C(_05869_),
    .X(_05921_));
 sky130_fd_sc_hd__and2_1 _12691_ (.A(_05920_),
    .B(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__o21ai_1 _12692_ (.A1(_05917_),
    .A2(_05918_),
    .B1(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__or3_1 _12693_ (.A(_05917_),
    .B(_05918_),
    .C(_05922_),
    .X(_05924_));
 sky130_fd_sc_hd__and2_1 _12694_ (.A(_05923_),
    .B(_05924_),
    .X(_05926_));
 sky130_fd_sc_hd__xnor2_1 _12695_ (.A(_05916_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__nand2_1 _12696_ (.A(_05915_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__or2_1 _12697_ (.A(_05915_),
    .B(_05927_),
    .X(_05929_));
 sky130_fd_sc_hd__nand2_1 _12698_ (.A(_05928_),
    .B(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__a21oi_2 _12699_ (.A1(_05852_),
    .A2(_05881_),
    .B1(_05850_),
    .Y(_05931_));
 sky130_fd_sc_hd__xnor2_1 _12700_ (.A(_05930_),
    .B(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__a21o_1 _12701_ (.A1(_05796_),
    .A2(_05812_),
    .B1(_05810_),
    .X(_05933_));
 sky130_fd_sc_hd__and2b_1 _12702_ (.A_N(_05853_),
    .B(_05880_),
    .X(_05934_));
 sky130_fd_sc_hd__nor2_1 _12703_ (.A(_05878_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__a2bb2o_2 _12704_ (.A1_N(_05251_),
    .A2_N(_05786_),
    .B1(_05787_),
    .B2(_05785_),
    .X(_05937_));
 sky130_fd_sc_hd__xor2_4 _12705_ (.A(_05775_),
    .B(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__nand2_1 _12706_ (.A(_05798_),
    .B(_05806_),
    .Y(_05939_));
 sky130_fd_sc_hd__or2b_1 _12707_ (.A(_05800_),
    .B_N(_05801_),
    .X(_05940_));
 sky130_fd_sc_hd__or2b_1 _12708_ (.A(_05601_),
    .B_N(_05856_),
    .X(_05941_));
 sky130_fd_sc_hd__o211a_1 _12709_ (.A1(_05857_),
    .A2(_05864_),
    .B1(_05862_),
    .C1(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__xnor2_1 _12710_ (.A(_05940_),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__a21o_1 _12711_ (.A1(_05803_),
    .A2(_05939_),
    .B1(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__nand3_1 _12712_ (.A(_05803_),
    .B(_05939_),
    .C(_05943_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_2 _12713_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__xor2_2 _12714_ (.A(_05938_),
    .B(_05946_),
    .X(_05948_));
 sky130_fd_sc_hd__xnor2_2 _12715_ (.A(_05935_),
    .B(_05948_),
    .Y(_05949_));
 sky130_fd_sc_hd__xor2_2 _12716_ (.A(_05933_),
    .B(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__xnor2_1 _12717_ (.A(_05932_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__and2b_1 _12718_ (.A_N(_05883_),
    .B(_05885_),
    .X(_05952_));
 sky130_fd_sc_hd__o21ba_1 _12719_ (.A1(_05815_),
    .A2(_05886_),
    .B1_N(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__xnor2_1 _12720_ (.A(_05951_),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__a21o_2 _12721_ (.A1(_05756_),
    .A2(_05759_),
    .B1(_05762_),
    .X(_05955_));
 sky130_fd_sc_hd__and2b_1 _12722_ (.A_N(_05813_),
    .B(_05770_),
    .X(_05956_));
 sky130_fd_sc_hd__a21o_1 _12723_ (.A1(_05768_),
    .A2(_05814_),
    .B1(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__a21boi_1 _12724_ (.A1(_05771_),
    .A2(_05779_),
    .B1_N(_05778_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ba_1 _12725_ (.A1(_05790_),
    .A2(_05793_),
    .B1_N(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__or3b_1 _12726_ (.A(_05790_),
    .B(_05793_),
    .C_N(_05959_),
    .X(_05961_));
 sky130_fd_sc_hd__and2b_2 _12727_ (.A_N(_05960_),
    .B(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__xor2_4 _12728_ (.A(_05757_),
    .B(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__xnor2_1 _12729_ (.A(_05957_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__xnor2_1 _12730_ (.A(_05955_),
    .B(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__xnor2_1 _12731_ (.A(_05954_),
    .B(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__nor2_1 _12732_ (.A(_05887_),
    .B(_05889_),
    .Y(_05967_));
 sky130_fd_sc_hd__a21oi_1 _12733_ (.A1(_05766_),
    .A2(_05890_),
    .B1(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__xnor2_1 _12734_ (.A(_05966_),
    .B(_05968_),
    .Y(_05970_));
 sky130_fd_sc_hd__or2b_1 _12735_ (.A(_05765_),
    .B_N(_05752_),
    .X(_05971_));
 sky130_fd_sc_hd__a21boi_1 _12736_ (.A1(_05754_),
    .A2(_05764_),
    .B1_N(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__xnor2_1 _12737_ (.A(_05970_),
    .B(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__a21oi_1 _12738_ (.A1(_05749_),
    .A2(_05895_),
    .B1(_05894_),
    .Y(_05974_));
 sky130_fd_sc_hd__or2_1 _12739_ (.A(_05973_),
    .B(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(_05973_),
    .B(_05974_),
    .Y(_05976_));
 sky130_fd_sc_hd__and2_1 _12741_ (.A(_05975_),
    .B(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__or2b_1 _12742_ (.A(_05898_),
    .B_N(_05897_),
    .X(_05978_));
 sky130_fd_sc_hd__and2b_1 _12743_ (.A_N(_05897_),
    .B(_05898_),
    .X(_05979_));
 sky130_fd_sc_hd__a21o_1 _12744_ (.A1(_05727_),
    .A2(_05978_),
    .B1(_05979_),
    .X(_05981_));
 sky130_fd_sc_hd__a31oi_2 _12745_ (.A1(_05730_),
    .A2(_05733_),
    .A3(_05899_),
    .B1(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__xnor2_1 _12746_ (.A(_05977_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__nand2_1 _12747_ (.A(net265),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__or2_1 _12748_ (.A(net265),
    .B(_05983_),
    .X(_05985_));
 sky130_fd_sc_hd__nand2_1 _12749_ (.A(_05984_),
    .B(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__inv_2 _12750_ (.A(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__or2_1 _12751_ (.A(net264),
    .B(_05900_),
    .X(_05988_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(net263),
    .A2(_05734_),
    .B1(_05900_),
    .B2(net264),
    .X(_05989_));
 sky130_fd_sc_hd__and3_1 _12753_ (.A(_05735_),
    .B(_05738_),
    .C(_05901_),
    .X(_05990_));
 sky130_fd_sc_hd__and3_1 _12754_ (.A(_05735_),
    .B(_05742_),
    .C(_05901_),
    .X(_05992_));
 sky130_fd_sc_hd__a221o_1 _12755_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_05990_),
    .B2(_05737_),
    .C1(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__or2_1 _12756_ (.A(_05987_),
    .B(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__nand2_1 _12757_ (.A(_05987_),
    .B(_05993_),
    .Y(_05995_));
 sky130_fd_sc_hd__and3_1 _12758_ (.A(_02174_),
    .B(_05994_),
    .C(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__clkbuf_1 _12759_ (.A(_05996_),
    .X(_00016_));
 sky130_fd_sc_hd__or2b_1 _12760_ (.A(_05913_),
    .B_N(_05910_),
    .X(_05997_));
 sky130_fd_sc_hd__o22a_1 _12761_ (.A1(_05821_),
    .A2(_05831_),
    .B1(_05907_),
    .B2(_05909_),
    .X(_05998_));
 sky130_fd_sc_hd__or2_2 _12762_ (.A(_05905_),
    .B(_05906_),
    .X(_05999_));
 sky130_fd_sc_hd__xnor2_1 _12763_ (.A(_05999_),
    .B(_05920_),
    .Y(_06000_));
 sky130_fd_sc_hd__xnor2_1 _12764_ (.A(_05998_),
    .B(_06000_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21oi_1 _12765_ (.A1(_05997_),
    .A2(_05928_),
    .B1(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__and3_1 _12766_ (.A(_05997_),
    .B(_05928_),
    .C(_06002_),
    .X(_06004_));
 sky130_fd_sc_hd__nor2_1 _12767_ (.A(_06003_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__o21a_1 _12768_ (.A1(_05938_),
    .A2(_05946_),
    .B1(_05944_),
    .X(_06006_));
 sky130_fd_sc_hd__or2b_1 _12769_ (.A(_05916_),
    .B_N(_05926_),
    .X(_06007_));
 sky130_fd_sc_hd__or2_2 _12770_ (.A(_05940_),
    .B(_05942_),
    .X(_06008_));
 sky130_fd_sc_hd__a21oi_1 _12771_ (.A1(_05923_),
    .A2(_06007_),
    .B1(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__and3_1 _12772_ (.A(_05923_),
    .B(_06007_),
    .C(_06008_),
    .X(_06010_));
 sky130_fd_sc_hd__nor2_1 _12773_ (.A(_06009_),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__xnor2_1 _12774_ (.A(_06006_),
    .B(_06011_),
    .Y(_06013_));
 sky130_fd_sc_hd__xnor2_1 _12775_ (.A(_06005_),
    .B(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _12776_ (.A(_05930_),
    .B(_05931_),
    .Y(_06015_));
 sky130_fd_sc_hd__nor2_1 _12777_ (.A(_05930_),
    .B(_05931_),
    .Y(_06016_));
 sky130_fd_sc_hd__a21oi_1 _12778_ (.A1(_06015_),
    .A2(_05950_),
    .B1(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__xnor2_1 _12779_ (.A(_06014_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__a21oi_4 _12780_ (.A1(_05757_),
    .A2(_05962_),
    .B1(_05960_),
    .Y(_06019_));
 sky130_fd_sc_hd__and3_2 _12781_ (.A(_05543_),
    .B(_05774_),
    .C(_05937_),
    .X(_06020_));
 sky130_fd_sc_hd__o21ai_1 _12782_ (.A1(_05878_),
    .A2(_05934_),
    .B1(_05948_),
    .Y(_06021_));
 sky130_fd_sc_hd__a21bo_1 _12783_ (.A1(_05933_),
    .A2(_05949_),
    .B1_N(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__xor2_1 _12784_ (.A(_06020_),
    .B(_06022_),
    .X(_06024_));
 sky130_fd_sc_hd__xnor2_1 _12785_ (.A(_06019_),
    .B(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__xor2_1 _12786_ (.A(_06018_),
    .B(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__and2b_1 _12787_ (.A_N(_05953_),
    .B(_05951_),
    .X(_06027_));
 sky130_fd_sc_hd__a21oi_1 _12788_ (.A1(_05954_),
    .A2(_05965_),
    .B1(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__or2_1 _12789_ (.A(_06026_),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__nand2_1 _12790_ (.A(_06026_),
    .B(_06028_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(_06029_),
    .B(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__and2b_1 _12792_ (.A_N(_05964_),
    .B(_05955_),
    .X(_06032_));
 sky130_fd_sc_hd__a21oi_1 _12793_ (.A1(_05957_),
    .A2(_05963_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__xnor2_1 _12794_ (.A(_06031_),
    .B(_06033_),
    .Y(_06035_));
 sky130_fd_sc_hd__or2_1 _12795_ (.A(_05966_),
    .B(_05968_),
    .X(_06036_));
 sky130_fd_sc_hd__o21a_1 _12796_ (.A1(_05970_),
    .A2(_05972_),
    .B1(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__nor2_1 _12797_ (.A(_06035_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__and2_1 _12798_ (.A(_06035_),
    .B(_06037_),
    .X(_06039_));
 sky130_fd_sc_hd__or2_1 _12799_ (.A(_06038_),
    .B(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__inv_2 _12800_ (.A(_05977_),
    .Y(_06041_));
 sky130_fd_sc_hd__o21a_1 _12801_ (.A1(_06041_),
    .A2(_05982_),
    .B1(_05975_),
    .X(_06042_));
 sky130_fd_sc_hd__xor2_1 _12802_ (.A(_06040_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__and2_1 _12803_ (.A(net266),
    .B(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__nor2_1 _12804_ (.A(net266),
    .B(_06043_),
    .Y(_06046_));
 sky130_fd_sc_hd__nor2_1 _12805_ (.A(_06044_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand2_1 _12806_ (.A(_05984_),
    .B(_05995_),
    .Y(_06048_));
 sky130_fd_sc_hd__a21o_1 _12807_ (.A1(_06047_),
    .A2(_06048_),
    .B1(_00166_),
    .X(_06049_));
 sky130_fd_sc_hd__o21ba_1 _12808_ (.A1(_06047_),
    .A2(_06048_),
    .B1_N(_06049_),
    .X(_00017_));
 sky130_fd_sc_hd__o21ba_1 _12809_ (.A1(_06040_),
    .A2(_06042_),
    .B1_N(_06038_),
    .X(_06050_));
 sky130_fd_sc_hd__a21o_1 _12810_ (.A1(_05999_),
    .A2(_05920_),
    .B1(_05998_),
    .X(_06051_));
 sky130_fd_sc_hd__o21ai_1 _12811_ (.A1(_05999_),
    .A2(_05920_),
    .B1(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__or2b_1 _12812_ (.A(_06019_),
    .B_N(_06024_),
    .X(_06053_));
 sky130_fd_sc_hd__a21bo_1 _12813_ (.A1(_06020_),
    .A2(_06022_),
    .B1_N(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__xnor2_1 _12814_ (.A(_06052_),
    .B(_06054_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21oi_1 _12815_ (.A1(_06005_),
    .A2(_06013_),
    .B1(_06003_),
    .Y(_06057_));
 sky130_fd_sc_hd__o21ai_1 _12816_ (.A1(_06031_),
    .A2(_06033_),
    .B1(_06029_),
    .Y(_06058_));
 sky130_fd_sc_hd__or2b_1 _12817_ (.A(_06018_),
    .B_N(_06025_),
    .X(_06059_));
 sky130_fd_sc_hd__o21a_1 _12818_ (.A1(_06014_),
    .A2(_06017_),
    .B1(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__xnor2_1 _12819_ (.A(_06058_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__and2b_1 _12820_ (.A_N(_06006_),
    .B(_06011_),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_1 _12821_ (.A(_06009_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_1 _12822_ (.A(_06061_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_1 _12823_ (.A(_06057_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__xnor2_2 _12824_ (.A(_06056_),
    .B(_06065_),
    .Y(_06067_));
 sky130_fd_sc_hd__xnor2_1 _12825_ (.A(_06050_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2_1 _12826_ (.A(net267),
    .B(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__nor2_1 _12827_ (.A(net267),
    .B(_06068_),
    .Y(_06070_));
 sky130_fd_sc_hd__nor2_1 _12828_ (.A(_06069_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__inv_2 _12829_ (.A(_05984_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21ba_1 _12830_ (.A1(_06072_),
    .A2(_06044_),
    .B1_N(_06046_),
    .X(_06073_));
 sky130_fd_sc_hd__a31o_1 _12831_ (.A1(_05987_),
    .A2(_05993_),
    .A3(_06047_),
    .B1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__or2_1 _12832_ (.A(_06071_),
    .B(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(_06071_),
    .B(_06074_),
    .Y(_06076_));
 sky130_fd_sc_hd__and3_1 _12834_ (.A(_02174_),
    .B(_06075_),
    .C(_06076_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _12835_ (.A(_06078_),
    .X(_00018_));
 sky130_fd_sc_hd__inv_2 _12836_ (.A(net268),
    .Y(_06079_));
 sky130_fd_sc_hd__a21oi_2 _12837_ (.A1(_06071_),
    .A2(_06074_),
    .B1(_06069_),
    .Y(_06080_));
 sky130_fd_sc_hd__nand2_1 _12838_ (.A(_06079_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__or2_1 _12839_ (.A(_06079_),
    .B(_06080_),
    .X(_06082_));
 sky130_fd_sc_hd__and3_1 _12840_ (.A(_02174_),
    .B(_06081_),
    .C(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _12841_ (.A(_06083_),
    .X(_00019_));
 sky130_fd_sc_hd__inv_2 _12842_ (.A(net270),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2_1 _12843_ (.A(_06084_),
    .B(_06082_),
    .Y(_06085_));
 sky130_fd_sc_hd__or2_1 _12844_ (.A(_06084_),
    .B(_06082_),
    .X(_06087_));
 sky130_fd_sc_hd__and3_1 _12845_ (.A(_02174_),
    .B(_06085_),
    .C(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _12846_ (.A(_06088_),
    .X(_00020_));
 sky130_fd_sc_hd__or2b_1 _12847_ (.A(net271),
    .B_N(_06087_),
    .X(_06089_));
 sky130_fd_sc_hd__or4b_4 _12848_ (.A(_06079_),
    .B(_06084_),
    .C(_06080_),
    .D_N(net271),
    .X(_06090_));
 sky130_fd_sc_hd__and3_1 _12849_ (.A(_02174_),
    .B(_06089_),
    .C(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _12850_ (.A(_06091_),
    .X(_00021_));
 sky130_fd_sc_hd__inv_2 _12851_ (.A(net272),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _12852_ (.A(_06092_),
    .B(_06090_),
    .Y(_06093_));
 sky130_fd_sc_hd__or2_1 _12853_ (.A(_06092_),
    .B(_06090_),
    .X(_06094_));
 sky130_fd_sc_hd__and3_1 _12854_ (.A(_02174_),
    .B(_06093_),
    .C(_06094_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _12855_ (.A(_06096_),
    .X(_00022_));
 sky130_fd_sc_hd__inv_2 _12856_ (.A(net273),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _12857_ (.A(_06097_),
    .B(_06094_),
    .Y(_06098_));
 sky130_fd_sc_hd__or3_4 _12858_ (.A(_06092_),
    .B(_06097_),
    .C(_06090_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_6 _12859_ (.A(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__and3_1 _12860_ (.A(_02174_),
    .B(_06098_),
    .C(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _12861_ (.A(_06101_),
    .X(_00023_));
 sky130_fd_sc_hd__inv_2 _12862_ (.A(net274),
    .Y(_06102_));
 sky130_fd_sc_hd__nor2_1 _12863_ (.A(_06102_),
    .B(_06100_),
    .Y(_06103_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_06102_),
    .B(_06100_),
    .Y(_06105_));
 sky130_fd_sc_hd__and3b_1 _12865_ (.A_N(_06103_),
    .B(_02174_),
    .C(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _12866_ (.A(_06106_),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _12867_ (.A(net274),
    .B(net275),
    .Y(_06107_));
 sky130_fd_sc_hd__o221a_1 _12868_ (.A1(net319),
    .A2(_06103_),
    .B1(_06107_),
    .B2(_06100_),
    .C1(_02185_),
    .X(_00025_));
 sky130_fd_sc_hd__nor2_1 _12869_ (.A(_06100_),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__inv_2 _12870_ (.A(net276),
    .Y(_06109_));
 sky130_fd_sc_hd__o31a_1 _12871_ (.A1(_06109_),
    .A2(_06100_),
    .A3(_06107_),
    .B1(_02185_),
    .X(_06110_));
 sky130_fd_sc_hd__o21a_1 _12872_ (.A1(net320),
    .A2(_06108_),
    .B1(_06110_),
    .X(_00026_));
 sky130_fd_sc_hd__o31ai_1 _12873_ (.A1(_06109_),
    .A2(_06100_),
    .A3(_06107_),
    .B1(net277),
    .Y(_06111_));
 sky130_fd_sc_hd__or4_4 _12874_ (.A(_06109_),
    .B(net277),
    .C(_06100_),
    .D(_06107_),
    .X(_06113_));
 sky130_fd_sc_hd__a21oi_2 _12875_ (.A1(_06111_),
    .A2(_06113_),
    .B1(_00166_),
    .Y(_00027_));
 sky130_fd_sc_hd__dfxtp_2 _12876_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00000_),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_2 _12877_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00001_),
    .Q(net269));
 sky130_fd_sc_hd__dfxtp_2 _12878_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00002_),
    .Q(net278));
 sky130_fd_sc_hd__dfxtp_1 _12879_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00003_),
    .Q(net279));
 sky130_fd_sc_hd__dfxtp_1 _12880_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00004_),
    .Q(net280));
 sky130_fd_sc_hd__dfxtp_1 _12881_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00005_),
    .Q(net281));
 sky130_fd_sc_hd__dfxtp_1 _12882_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00006_),
    .Q(net282));
 sky130_fd_sc_hd__dfxtp_1 _12883_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00007_),
    .Q(net283));
 sky130_fd_sc_hd__dfxtp_1 _12884_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00008_),
    .Q(net284));
 sky130_fd_sc_hd__dfxtp_1 _12885_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00009_),
    .Q(net285));
 sky130_fd_sc_hd__dfxtp_1 _12886_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00010_),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_1 _12887_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00011_),
    .Q(net260));
 sky130_fd_sc_hd__dfxtp_1 _12888_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00012_),
    .Q(net261));
 sky130_fd_sc_hd__dfxtp_1 _12889_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00013_),
    .Q(net262));
 sky130_fd_sc_hd__dfxtp_1 _12890_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00014_),
    .Q(net263));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00015_),
    .Q(net264));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00016_),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00017_),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00018_),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00019_),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00020_),
    .Q(net270));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00021_),
    .Q(net271));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00022_),
    .Q(net272));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00023_),
    .Q(net273));
 sky130_fd_sc_hd__dfxtp_1 _12900_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00024_),
    .Q(net274));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00025_),
    .Q(net275));
 sky130_fd_sc_hd__dfxtp_1 _12902_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00026_),
    .Q(net276));
 sky130_fd_sc_hd__dfxtp_1 _12903_ (.CLK(clknet_1_1__leaf_clk),
    .D(_00027_),
    .Q(net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net275),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net276),
    .X(net320));
 sky130_fd_sc_hd__buf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(data_in[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(data_in[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(data_in[190]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(data_in[191]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(data_in[192]),
    .X(net103));
 sky130_fd_sc_hd__buf_4 input104 (.A(data_in[193]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(data_in[194]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(data_in[195]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(data_in[196]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(data_in[197]),
    .X(net108));
 sky130_fd_sc_hd__buf_4 input109 (.A(data_in[198]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(data_in[109]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(data_in[199]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(data_in[19]),
    .X(net111));
 sky130_fd_sc_hd__buf_4 input112 (.A(data_in[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(data_in[200]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(data_in[201]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(data_in[202]),
    .X(net115));
 sky130_fd_sc_hd__buf_4 input116 (.A(data_in[203]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(data_in[204]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 input118 (.A(data_in[205]),
    .X(net118));
 sky130_fd_sc_hd__buf_4 input119 (.A(data_in[206]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(data_in[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input120 (.A(data_in[207]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(data_in[208]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(data_in[209]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(data_in[20]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 input124 (.A(data_in[210]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 input125 (.A(data_in[211]),
    .X(net125));
 sky130_fd_sc_hd__buf_2 input126 (.A(data_in[212]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input127 (.A(data_in[213]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(data_in[214]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(data_in[215]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(data_in[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input130 (.A(data_in[216]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(data_in[217]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(data_in[218]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(data_in[219]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(data_in[21]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(data_in[220]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(data_in[221]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(data_in[222]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(data_in[223]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(data_in[224]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input14 (.A(data_in[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input140 (.A(data_in[225]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(data_in[226]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(data_in[227]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(data_in[228]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(data_in[229]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 input145 (.A(data_in[22]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(data_in[230]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(data_in[231]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(data_in[232]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(data_in[233]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(data_in[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input150 (.A(data_in[234]),
    .X(net150));
 sky130_fd_sc_hd__buf_2 input151 (.A(data_in[235]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(data_in[236]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(data_in[237]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(data_in[238]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(data_in[239]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(data_in[23]),
    .X(net156));
 sky130_fd_sc_hd__buf_2 input157 (.A(data_in[240]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(data_in[241]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(data_in[242]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(data_in[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input160 (.A(data_in[243]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(data_in[244]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(data_in[245]),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(data_in[246]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(data_in[247]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(data_in[248]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 input166 (.A(data_in[249]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(data_in[24]),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(data_in[250]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(data_in[251]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(data_in[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input170 (.A(data_in[252]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(data_in[253]),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(data_in[254]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 input173 (.A(data_in[255]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 input174 (.A(data_in[25]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 input175 (.A(data_in[26]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 input176 (.A(data_in[27]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 input177 (.A(data_in[28]),
    .X(net177));
 sky130_fd_sc_hd__buf_4 input178 (.A(data_in[29]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(data_in[2]),
    .X(net179));
 sky130_fd_sc_hd__buf_4 input18 (.A(data_in[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input180 (.A(data_in[30]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(data_in[31]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 input182 (.A(data_in[32]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 input183 (.A(data_in[33]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 input184 (.A(data_in[34]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(data_in[35]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 input186 (.A(data_in[36]),
    .X(net186));
 sky130_fd_sc_hd__buf_2 input187 (.A(data_in[37]),
    .X(net187));
 sky130_fd_sc_hd__buf_4 input188 (.A(data_in[38]),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(data_in[39]),
    .X(net189));
 sky130_fd_sc_hd__buf_4 input19 (.A(data_in[116]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(data_in[3]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 input191 (.A(data_in[40]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 input192 (.A(data_in[41]),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input193 (.A(data_in[42]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(data_in[43]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(data_in[44]),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(data_in[45]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input197 (.A(data_in[46]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(data_in[47]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(data_in[48]),
    .X(net199));
 sky130_fd_sc_hd__buf_2 input2 (.A(data_in[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input20 (.A(data_in[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input200 (.A(data_in[49]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(data_in[4]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(data_in[50]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(data_in[51]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 input204 (.A(data_in[52]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 input205 (.A(data_in[53]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(data_in[54]),
    .X(net206));
 sky130_fd_sc_hd__buf_2 input207 (.A(data_in[55]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(data_in[56]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 input209 (.A(data_in[57]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(data_in[118]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input210 (.A(data_in[58]),
    .X(net210));
 sky130_fd_sc_hd__buf_2 input211 (.A(data_in[59]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(data_in[5]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(data_in[60]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(data_in[61]),
    .X(net214));
 sky130_fd_sc_hd__buf_2 input215 (.A(data_in[62]),
    .X(net215));
 sky130_fd_sc_hd__buf_4 input216 (.A(data_in[63]),
    .X(net216));
 sky130_fd_sc_hd__buf_2 input217 (.A(data_in[64]),
    .X(net217));
 sky130_fd_sc_hd__buf_2 input218 (.A(data_in[65]),
    .X(net218));
 sky130_fd_sc_hd__buf_2 input219 (.A(data_in[66]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(data_in[119]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input220 (.A(data_in[67]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 input221 (.A(data_in[68]),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(data_in[69]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(data_in[6]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(data_in[70]),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(data_in[71]),
    .X(net225));
 sky130_fd_sc_hd__buf_2 input226 (.A(data_in[72]),
    .X(net226));
 sky130_fd_sc_hd__buf_2 input227 (.A(data_in[73]),
    .X(net227));
 sky130_fd_sc_hd__buf_4 input228 (.A(data_in[74]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 input229 (.A(data_in[75]),
    .X(net229));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(data_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(data_in[76]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input231 (.A(data_in[77]),
    .X(net231));
 sky130_fd_sc_hd__buf_2 input232 (.A(data_in[78]),
    .X(net232));
 sky130_fd_sc_hd__buf_2 input233 (.A(data_in[79]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(data_in[7]),
    .X(net234));
 sky130_fd_sc_hd__buf_2 input235 (.A(data_in[80]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 input236 (.A(data_in[81]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 input237 (.A(data_in[82]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 input238 (.A(data_in[83]),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input239 (.A(data_in[84]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(data_in[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input240 (.A(data_in[85]),
    .X(net240));
 sky130_fd_sc_hd__buf_2 input241 (.A(data_in[86]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(data_in[87]),
    .X(net242));
 sky130_fd_sc_hd__buf_2 input243 (.A(data_in[88]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 input244 (.A(data_in[89]),
    .X(net244));
 sky130_fd_sc_hd__buf_4 input245 (.A(data_in[8]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 input246 (.A(data_in[90]),
    .X(net246));
 sky130_fd_sc_hd__buf_2 input247 (.A(data_in[91]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 input248 (.A(data_in[92]),
    .X(net248));
 sky130_fd_sc_hd__buf_2 input249 (.A(data_in[93]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(data_in[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input250 (.A(data_in[94]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 input251 (.A(data_in[95]),
    .X(net251));
 sky130_fd_sc_hd__buf_2 input252 (.A(data_in[96]),
    .X(net252));
 sky130_fd_sc_hd__dlymetal6s2s_1 input253 (.A(data_in[97]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 input254 (.A(data_in[98]),
    .X(net254));
 sky130_fd_sc_hd__buf_2 input255 (.A(data_in[99]),
    .X(net255));
 sky130_fd_sc_hd__buf_6 input256 (.A(data_in[9]),
    .X(net256));
 sky130_fd_sc_hd__buf_4 input257 (.A(reset),
    .X(net257));
 sky130_fd_sc_hd__buf_4 input26 (.A(data_in[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(data_in[123]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(data_in[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(data_in[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(data_in[101]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(data_in[126]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(data_in[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(data_in[128]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(data_in[129]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(data_in[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(data_in[130]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(data_in[131]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(data_in[132]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(data_in[133]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(data_in[134]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(data_in[102]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(data_in[135]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(data_in[136]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(data_in[137]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(data_in[138]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(data_in[139]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(data_in[13]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(data_in[140]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(data_in[141]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(data_in[142]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(data_in[143]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(data_in[103]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(data_in[144]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(data_in[145]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(data_in[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(data_in[147]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(data_in[148]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(data_in[149]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(data_in[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(data_in[150]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(data_in[151]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(data_in[152]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(data_in[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input60 (.A(data_in[153]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(data_in[154]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(data_in[155]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(data_in[156]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(data_in[157]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(data_in[158]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(data_in[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(data_in[15]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(data_in[160]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(data_in[161]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(data_in[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input70 (.A(data_in[162]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(data_in[163]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(data_in[164]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(data_in[165]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 input74 (.A(data_in[166]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(data_in[167]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(data_in[168]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(data_in[169]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(data_in[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(data_in[170]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(data_in[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input80 (.A(data_in[171]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(data_in[172]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(data_in[173]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(data_in[174]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(data_in[175]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(data_in[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(data_in[177]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(data_in[178]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(data_in[179]),
    .X(net88));
 sky130_fd_sc_hd__buf_4 input89 (.A(data_in[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(data_in[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(data_in[180]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(data_in[181]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(data_in[182]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(data_in[183]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(data_in[184]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(data_in[185]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(data_in[186]),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input97 (.A(data_in[187]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(data_in[188]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(data_in[189]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 max_cap1 (.A(_01115_),
    .X(net318));
 sky130_fd_sc_hd__buf_1 max_cap286 (.A(_01714_),
    .X(net286));
 sky130_fd_sc_hd__buf_1 max_cap287 (.A(_01115_),
    .X(net287));
 sky130_fd_sc_hd__buf_1 max_cap288 (.A(net322),
    .X(net288));
 sky130_fd_sc_hd__buf_1 max_cap289 (.A(_00801_),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 max_cap290 (.A(_01111_),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 max_cap291 (.A(_01107_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 max_cap292 (.A(_00736_),
    .X(net292));
 sky130_fd_sc_hd__buf_1 max_cap293 (.A(_02579_),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 max_cap294 (.A(_01103_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 max_cap295 (.A(_00792_),
    .X(net295));
 sky130_fd_sc_hd__buf_1 max_cap296 (.A(_00412_),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 max_cap297 (.A(_00137_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 max_cap298 (.A(_00866_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 max_cap299 (.A(_00573_),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(_00149_),
    .X(net322));
 sky130_fd_sc_hd__buf_1 max_cap300 (.A(net324),
    .X(net300));
 sky130_fd_sc_hd__buf_1 max_cap301 (.A(_01095_),
    .X(net301));
 sky130_fd_sc_hd__buf_1 max_cap302 (.A(_00569_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 max_cap304 (.A(_02233_),
    .X(net304));
 sky130_fd_sc_hd__buf_1 max_cap305 (.A(_02091_),
    .X(net305));
 sky130_fd_sc_hd__buf_1 max_cap306 (.A(_01091_),
    .X(net306));
 sky130_fd_sc_hd__buf_1 max_cap308 (.A(_06269_),
    .X(net308));
 sky130_fd_sc_hd__buf_1 max_cap4 (.A(_01103_),
    .X(net323));
 sky130_fd_sc_hd__buf_1 max_cap5 (.A(_01095_),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .X(data_out[10]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(data_out[11]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(data_out[12]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(data_out[13]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(data_out[14]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(data_out[15]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .X(data_out[16]));
 sky130_fd_sc_hd__clkbuf_4 output266 (.A(net266),
    .X(data_out[17]));
 sky130_fd_sc_hd__clkbuf_4 output267 (.A(net267),
    .X(data_out[18]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .X(data_out[19]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .X(data_out[20]));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net271),
    .X(data_out[21]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .X(data_out[22]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .X(data_out[23]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .X(data_out[24]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(data_out[25]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(data_out[26]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .X(data_out[27]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(data_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(data_out[9]));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer1 (.A(_00581_),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(_00584_),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(_01688_),
    .X(net310));
 sky130_fd_sc_hd__buf_1 rebuffer3 (.A(_01688_),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(net325),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(_00600_),
    .X(net313));
 sky130_fd_sc_hd__buf_1 rebuffer6 (.A(_00579_),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(_00117_),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(_00116_),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(_00119_),
    .X(net317));
 sky130_fd_sc_hd__buf_1 wire2 (.A(_01111_),
    .X(net321));
 sky130_fd_sc_hd__buf_1 wire303 (.A(_00181_),
    .X(net303));
 sky130_fd_sc_hd__buf_1 wire307 (.A(_00069_),
    .X(net307));
endmodule

