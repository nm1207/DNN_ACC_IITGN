* NGSPICE file created from mac.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt mac VGND VPWR clk data_in[0] data_in[100] data_in[101] data_in[102] data_in[103]
+ data_in[104] data_in[105] data_in[106] data_in[107] data_in[108] data_in[109] data_in[10]
+ data_in[110] data_in[111] data_in[112] data_in[113] data_in[114] data_in[115] data_in[116]
+ data_in[117] data_in[118] data_in[119] data_in[11] data_in[120] data_in[121] data_in[122]
+ data_in[123] data_in[124] data_in[125] data_in[126] data_in[127] data_in[128] data_in[129]
+ data_in[12] data_in[130] data_in[131] data_in[132] data_in[133] data_in[134] data_in[135]
+ data_in[136] data_in[137] data_in[138] data_in[139] data_in[13] data_in[140] data_in[141]
+ data_in[142] data_in[143] data_in[144] data_in[145] data_in[146] data_in[147] data_in[148]
+ data_in[149] data_in[14] data_in[150] data_in[151] data_in[152] data_in[153] data_in[154]
+ data_in[155] data_in[156] data_in[157] data_in[158] data_in[159] data_in[15] data_in[160]
+ data_in[161] data_in[162] data_in[163] data_in[164] data_in[165] data_in[166] data_in[167]
+ data_in[168] data_in[169] data_in[16] data_in[170] data_in[171] data_in[172] data_in[173]
+ data_in[174] data_in[175] data_in[176] data_in[177] data_in[178] data_in[179] data_in[17]
+ data_in[180] data_in[181] data_in[182] data_in[183] data_in[184] data_in[185] data_in[186]
+ data_in[187] data_in[188] data_in[189] data_in[18] data_in[190] data_in[191] data_in[192]
+ data_in[193] data_in[194] data_in[195] data_in[196] data_in[197] data_in[198] data_in[199]
+ data_in[19] data_in[1] data_in[200] data_in[201] data_in[202] data_in[203] data_in[204]
+ data_in[205] data_in[206] data_in[207] data_in[208] data_in[209] data_in[20] data_in[210]
+ data_in[211] data_in[212] data_in[213] data_in[214] data_in[215] data_in[216] data_in[217]
+ data_in[218] data_in[219] data_in[21] data_in[220] data_in[221] data_in[222] data_in[223]
+ data_in[224] data_in[225] data_in[226] data_in[227] data_in[228] data_in[229] data_in[22]
+ data_in[230] data_in[231] data_in[232] data_in[233] data_in[234] data_in[235] data_in[236]
+ data_in[237] data_in[238] data_in[239] data_in[23] data_in[240] data_in[241] data_in[242]
+ data_in[243] data_in[244] data_in[245] data_in[246] data_in[247] data_in[248] data_in[249]
+ data_in[24] data_in[250] data_in[251] data_in[252] data_in[253] data_in[254] data_in[255]
+ data_in[25] data_in[26] data_in[27] data_in[28] data_in[29] data_in[2] data_in[30]
+ data_in[31] data_in[32] data_in[33] data_in[34] data_in[35] data_in[36] data_in[37]
+ data_in[38] data_in[39] data_in[3] data_in[40] data_in[41] data_in[42] data_in[43]
+ data_in[44] data_in[45] data_in[46] data_in[47] data_in[48] data_in[49] data_in[4]
+ data_in[50] data_in[51] data_in[52] data_in[53] data_in[54] data_in[55] data_in[56]
+ data_in[57] data_in[58] data_in[59] data_in[5] data_in[60] data_in[61] data_in[62]
+ data_in[63] data_in[64] data_in[65] data_in[66] data_in[67] data_in[68] data_in[69]
+ data_in[6] data_in[70] data_in[71] data_in[72] data_in[73] data_in[74] data_in[75]
+ data_in[76] data_in[77] data_in[78] data_in[79] data_in[7] data_in[80] data_in[81]
+ data_in[82] data_in[83] data_in[84] data_in[85] data_in[86] data_in[87] data_in[88]
+ data_in[89] data_in[8] data_in[90] data_in[91] data_in[92] data_in[93] data_in[94]
+ data_in[95] data_in[96] data_in[97] data_in[98] data_in[99] data_in[9] data_out[0]
+ data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16]
+ data_out[17] data_out[18] data_out[19] data_out[1] data_out[20] data_out[21] data_out[22]
+ data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[2] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] reset
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09671_ _02606_ _02608_ _02586_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__o21a_1
X_06883_ _06195_ _06196_ _04029_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__o21ai_2
X_08622_ _01521_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08553_ _00885_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08484_ net240 VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07504_ _00385_ _06433_ _00405_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07435_ _00335_ _00336_ _06404_ _06406_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07366_ net308 VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__inv_2
X_09105_ net247 _00834_ _00366_ net238 VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__a22o_1
X_07297_ net90 VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09036_ _01299_ _01301_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09938_ net198 VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09869_ _02826_ _02827_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__and2b_1
X_11900_ _01666_ _03006_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__nand2_2
X_12880_ clknet_1_0__leaf_clk _00004_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dfxtp_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _00937_ _02799_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__and3_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11762_ _04894_ _04903_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _04815_ _04400_ _04826_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__or3_1
X_10713_ net19 _00706_ _00647_ _01181_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand4_1
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10644_ _03675_ _03677_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__xor2_2
X_10575_ _03004_ _03005_ _03007_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer7 _00117_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12314_ _05199_ _05232_ _05508_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12245_ _01562_ _02239_ _02904_ _01584_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12176_ _05355_ _05357_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__and3_1
X_11127_ _03600_ _03652_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a21bo_2
X_11058_ _04130_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__xor2_2
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10009_ net37 net46 _01051_ net36 VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07220_ _02811_ _00107_ _00121_ _00122_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07151_ _05158_ _00053_ _00054_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07082_ _06367_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07984_ _02569_ _00879_ _00883_ _00884_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09723_ _02055_ _02102_ _02101_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__a21bo_2
X_06935_ _06247_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09654_ net155 VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__clkbuf_4
X_06866_ _06178_ _04150_ _02394_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08605_ _01503_ _01504_ _01497_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__a21o_1
X_06797_ _06066_ _06095_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__xor2_2
X_09585_ _02513_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__nand2_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _02580_ _01434_ _01435_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08467_ net235 _01367_ _01365_ net208 VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_135_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08398_ _01292_ _01294_ _01297_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__o211ai_2
X_07418_ _00318_ _00319_ _06322_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07349_ _06263_ _00249_ _00251_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10360_ _06368_ net4 net5 _05882_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09019_ _06362_ _06304_ _01324_ _01325_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__and4_1
X_10291_ _03288_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12030_ _05184_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__xor2_4
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12863_ _06102_ _06100_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__nor2_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12794_ _06031_ _06033_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__xnor2_1
X_11814_ _04946_ _04960_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__xnor2_2
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _04883_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11676_ _04808_ _04809_ _04355_ _04363_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10627_ _02947_ _03040_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10558_ _03578_ _03581_ _03582_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12228_ _01653_ _04154_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nand2_1
X_10489_ _02873_ _02875_ _03506_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__a211oi_4
X_12159_ _05322_ _05338_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06720_ _05246_ _05257_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06651_ _04490_ _04501_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__nor2_1
X_09370_ _02278_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06582_ _03732_ _02569_ _03743_ _02580_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08321_ _01216_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08252_ _00172_ _00622_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__nand2_1
X_07203_ net36 VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08183_ _01081_ _01082_ _01083_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07134_ _06434_ _06435_ _00036_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07065_ _05893_ _05947_ _05936_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput264 net264 VGND VGND VPWR VPWR data_out[15] sky130_fd_sc_hd__clkbuf_4
Xoutput275 net275 VGND VGND VPWR VPWR data_out[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07967_ _00430_ _00451_ _00868_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__o21ai_2
X_09706_ _02609_ _02610_ _02645_ _02647_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__a2bb2o_1
X_06918_ _04490_ _06132_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__and3_1
X_07898_ _00797_ _00798_ _00414_ _00417_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a211oi_1
X_09637_ _01886_ _01888_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06849_ _06150_ _06163_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09568_ _01834_ _01842_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__or2_1
X_08519_ _00857_ _00859_ _00856_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__a21o_1
X_11530_ _04647_ _04650_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09499_ net169 net161 _00171_ _01777_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__nand4_1
XFILLER_0_37_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire303 _00181_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11461_ _04065_ _04067_ _04066_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11392_ _04026_ _04036_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__a21o_1
X_10412_ _02751_ _02783_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10343_ net2 net11 net13 net255 VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10274_ _03262_ _03269_ _03270_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12013_ _04842_ _04886_ _04883_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap5 _01095_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12846_ _06088_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12777_ _05930_ _05931_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__nor2_1
X_11728_ _04865_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _04768_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08870_ _01179_ _01197_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07821_ _00721_ _00722_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__xnor2_1
X_07752_ _00256_ _00653_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06703_ _03337_ _02712_ _03348_ _02723_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__and4_1
X_07683_ _00583_ _00584_ _00418_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__o21a_1
X_09422_ _01655_ _02336_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__xnor2_2
X_06634_ _04303_ _02218_ _04314_ _02229_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a22o_2
XFILLER_0_94_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _02200_ _02259_ _02260_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__nor3_1
X_08304_ _06138_ _00250_ _01202_ _01203_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__nand4_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06565_ _02646_ _03535_ _03557_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06496_ net41 VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09284_ _02159_ _02183_ _02184_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08235_ _01135_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08166_ net38 VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07117_ _06429_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08097_ _00996_ _00997_ _00484_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a21oi_1
X_07048_ _06361_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08999_ _01341_ _01343_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__and2b_1
X_10961_ _03442_ _03444_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nand2_2
X_12700_ _05930_ _05931_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__xnor2_1
X_10892_ _06375_ _02019_ _03947_ _03948_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nand4_2
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12631_ _05601_ _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12562_ _05771_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__xor2_1
X_11513_ _04604_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12493_ _05453_ _05456_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11444_ _04047_ _04048_ _04050_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__or3_2
XFILLER_0_61_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11375_ _03966_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10326_ _03327_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nand2_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10257_ _02645_ _02648_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__nand2_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10188_ _03175_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12829_ _05984_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08020_ _05389_ _05444_ _06437_ _06416_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09971_ _02235_ _02249_ _02248_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__a21boi_2
X_08922_ _06261_ net28 _01820_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08853_ _01751_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08784_ _01682_ _01683_ _01648_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__a21bo_1
X_07804_ net20 VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__buf_2
X_07735_ _00613_ _00636_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__xnor2_2
X_07666_ _00542_ _00567_ _00568_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__nor3_1
X_09405_ _02315_ _02316_ _02310_ _02311_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__a211o_1
X_06617_ net149 VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__clkbuf_4
X_07597_ _00488_ _00499_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09336_ net193 _01002_ _02238_ _02241_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__nand4_2
X_06548_ net89 VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09267_ _02164_ _02165_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08218_ _01117_ _01118_ _00637_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__a21oi_1
X_06479_ _02602_ _02613_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09198_ _02095_ _02096_ _01513_ _01515_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08149_ net47 VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__buf_4
X_11160_ _04243_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11091_ _01068_ _01051_ _01653_ _00530_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a22oi_1
X_10111_ _02454_ _02483_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10042_ _03016_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__xor2_4
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11993_ _04273_ _04740_ _04745_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__a21o_1
X_10944_ _04004_ _04006_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__xor2_2
X_10875_ _03328_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__xor2_4
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12614_ _05666_ _05673_ _05671_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a21o_2
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12545_ _05755_ _05760_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12476_ _05686_ _05687_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__nand2_2
X_11427_ _00937_ _01488_ _02799_ _00421_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ _00357_ _02019_ _04460_ _04461_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10309_ _03308_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__nor2_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _03878_ _03901_ _04385_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a21o_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07520_ _03579_ _02668_ _06410_ _00421_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07451_ _00352_ _00353_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07382_ _06145_ _06249_ _00283_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09121_ _03820_ _05914_ _00821_ net13 VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__nand4_2
XFILLER_0_57_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09052_ _01949_ _01950_ _01937_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08003_ _00806_ _00903_ _00904_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__nor3_2
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap296 _00412_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09954_ _02917_ _02918_ _02919_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__a21o_1
X_08905_ _01259_ _01260_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__or2b_1
X_09885_ _02829_ _02843_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__or3_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _01189_ _01191_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08767_ _02789_ _03106_ _01666_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__nand4_2
X_08698_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__or2b_1
X_07718_ _00273_ _00275_ _00619_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__or3_1
X_07649_ net256 net190 net201 net245 VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10660_ _03693_ _03694_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand2_2
XFILLER_0_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09319_ _05115_ _01567_ _02221_ _02222_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__nand4_2
XFILLER_0_63_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10591_ _03095_ _04939_ _01652_ _03006_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _05524_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__xnor2_1
X_12261_ _05431_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__xor2_4
XFILLER_0_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11212_ _03751_ _03759_ _03760_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a31oi_2
X_12192_ _05374_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11143_ _03316_ _03670_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__a21oi_4
Xinput120 data_in[207] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
X_11074_ _04148_ _04149_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__xor2_2
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput142 data_in[227] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
Xinput131 data_in[217] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput153 data_in[237] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
X_10025_ _02996_ _02997_ _02981_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a21o_1
Xinput175 data_in[26] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_4
Xinput164 data_in[247] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
Xinput186 data_in[36] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_4
Xinput197 data_in[46] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11976_ _05138_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__nand2_1
X_10927_ net55 net64 net57 net63 VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10858_ _03848_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__xnor2_2
X_10789_ _03814_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__xnor2_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12528_ _05735_ _05743_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12459_ _02239_ _02904_ _05667_ _05413_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06951_ _04435_ _02207_ _06142_ _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__nand4_2
X_09670_ _02586_ _02606_ _02608_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08621_ net113 net114 net108 net109 VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__and4_1
X_06882_ _04029_ _06195_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__or3_2
X_08552_ _01447_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08483_ _01382_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__and2_1
X_07503_ _00385_ _06433_ _00405_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07434_ _06404_ _06406_ _00335_ _00336_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07365_ _00267_ _04479_ _06247_ _06248_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__or4_1
X_09104_ net238 net247 _00366_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__and3_1
X_07296_ _06282_ _06287_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__and2b_1
X_09035_ _01932_ _01933_ _01333_ _01335_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09937_ _02901_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nor2_1
X_09868_ _02824_ _02825_ _02819_ _02820_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a211o_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _02126_ _02156_ _02155_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__a21boi_2
X_08819_ net282 _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__and2_1
X_11830_ _00421_ _01488_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__nand2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11761_ _04901_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10712_ net20 net29 net30 net19 VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a22o_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _04815_ _04400_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10643_ _02451_ _03054_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__a21oi_2
X_10574_ _02994_ _02996_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__or2b_2
XFILLER_0_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer8 _00116_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12313_ _05231_ _05229_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12244_ _05033_ _05035_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ _04988_ _04989_ _04987_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11126_ _03651_ _03649_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11057_ _03553_ _03561_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10008_ _01655_ _02335_ _02334_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__a21o_1
X_11959_ _04709_ _04712_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07150_ _00051_ _00052_ _05126_ _05147_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07081_ _06382_ _06394_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07983_ _02569_ _00879_ _00883_ _00884_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__nand4_2
X_09722_ _02453_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__xor2_4
X_06934_ _06244_ _06245_ _06246_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__nor3_1
X_09653_ _00749_ _02588_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__a21bo_1
X_06865_ _04128_ _04139_ _06178_ _02383_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__a22o_1
X_09584_ _02511_ _02512_ _02495_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__a21o_1
X_08604_ _01497_ _01503_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__nand3_2
X_08535_ _03732_ _05750_ _00397_ _00872_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__nand4_2
X_06796_ _02448_ _06086_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ net250 VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08397_ _06177_ _01293_ _01295_ _01296_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__nand4_4
X_07417_ _06322_ _00318_ _00319_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07348_ net15 _00250_ _00247_ _00248_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07279_ _06148_ _06251_ _00180_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__o21a_1
X_09018_ _04106_ _06173_ _00343_ _00810_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__and4_1
X_10290_ _06362_ _02626_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12862_ net274 VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__inv_2
X_11813_ _04952_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ _05957_ _05963_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a21oi_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11744_ _04880_ _04882_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11675_ _04354_ _04361_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__and2_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _03039_ _03037_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10557_ _03578_ _03581_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10488_ _03504_ _03505_ _02920_ _02923_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12227_ _04679_ _04681_ _05087_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__o21ba_1
X_12158_ _05322_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nor2_1
X_11109_ _04186_ _04187_ _03022_ _03639_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__a211o_1
X_12089_ _05240_ _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__xor2_2
X_06650_ _02251_ _04424_ _04457_ _04479_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06581_ net60 VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__buf_2
X_08320_ _01219_ _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08251_ _01150_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07202_ _02811_ _04906_ _04983_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08182_ _01081_ _01082_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ _06434_ _06435_ _00036_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07064_ _06372_ _06377_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput265 net265 VGND VGND VPWR VPWR data_out[16] sky130_fd_sc_hd__clkbuf_4
Xoutput276 net276 VGND VGND VPWR VPWR data_out[26] sky130_fd_sc_hd__clkbuf_4
X_07966_ _00449_ _00450_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__or2b_1
X_09705_ _02609_ _02610_ _02645_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06917_ _06229_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__nor2_1
X_09636_ _02543_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__xor2_4
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07897_ _00414_ _00417_ _00797_ _00798_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__o211a_1
X_06848_ _06161_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__xnor2_1
X_06779_ net254 VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09567_ _01840_ _01841_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__nand2_1
X_08518_ _01416_ _01417_ _01405_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__a21o_1
X_09498_ net161 net170 net162 net169 VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__a22o_1
X_08449_ _01347_ _01348_ _00790_ net295 VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11460_ _00985_ _01524_ _04571_ _04572_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10411_ _03387_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__xnor2_2
X_11391_ _04027_ _04035_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10342_ _02708_ _02710_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10273_ _03266_ _03267_ _03268_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12012_ _05176_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__nor2_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _02174_ _06085_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and3_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12776_ _05930_ _05931_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__nand2_1
X_11727_ _00757_ _01365_ _02626_ _01986_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__nand4_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ _04769_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10609_ _03638_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11589_ _03739_ _04228_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07820_ _04424_ _06159_ _06134_ _06284_ _00230_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__a41o_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07751_ _00651_ _00652_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__and2_1
X_06702_ _04730_ _05060_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07682_ _00418_ _00583_ net325 VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__nor3_2
X_09421_ _02334_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06633_ net131 VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__clkbuf_4
X_09352_ _02257_ _02258_ _02201_ _01626_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__a211oi_1
X_06564_ _03524_ _02635_ _03546_ _02646_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__a22o_1
X_08303_ _06138_ _00250_ _01202_ _01203_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06495_ net1 VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09283_ _02181_ _02182_ _02160_ _02161_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o211ai_2
X_08234_ _00613_ _00635_ _00634_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__o21bai_1
X_08165_ _01049_ _01050_ _01064_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07116_ _06421_ _06422_ _06428_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08096_ _00484_ _00996_ _00997_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__and3_1
X_07047_ net203 VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08998_ _01284_ _01345_ _01346_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nor3_2
X_07949_ _03798_ _00357_ _00850_ _02470_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__a22o_1
X_10960_ _03567_ _03521_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__and2b_1
X_10891_ _06375_ net14 _03947_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a22o_1
X_09619_ net125 _00665_ _02551_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__a22o_1
X_12630_ _02694_ _01367_ _02695_ _01987_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__and4_1
XFILLER_0_65_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12561_ _05778_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11512_ _04618_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12492_ _05679_ _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11443_ _04553_ _04554_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__or2_4
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11374_ _04475_ _04478_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__xnor2_2
X_10325_ net237 net238 net250 net251 VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__nand4_4
XFILLER_0_21_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10256_ _02687_ _02748_ _03251_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__o21a_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ _03173_ _03174_ net88 net101 VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12828_ _06069_ _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12759_ _05996_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09970_ _02926_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__xor2_2
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08921_ net26 net27 net19 net20 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08852_ _01155_ _01158_ _01154_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__o21ba_1
X_07803_ _04292_ net85 _00238_ _00703_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__nand4_2
X_08783_ _01648_ _01682_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_79_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07734_ _00634_ _00635_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07665_ _00563_ _00564_ _00566_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__a21oi_2
X_06616_ net140 VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__buf_2
X_09404_ _02310_ _02311_ _02315_ _02316_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07596_ _00496_ _00498_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09335_ _05093_ _01002_ _02238_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__a22o_1
X_06547_ _03337_ _02712_ _03348_ _02723_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nand4_1
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09266_ net78 net181 net110 net113 VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__a22o_1
X_06478_ _02558_ _02591_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08217_ _00637_ _01117_ _01118_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09197_ _01513_ _01515_ _02095_ _02096_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08148_ _00531_ _00538_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08079_ _00979_ _00980_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11090_ _03621_ _03625_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__and2_1
X_10110_ _02482_ _02455_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__or2b_1
X_10041_ _00549_ _01072_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11992_ _04790_ _04768_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__or2b_1
X_10943_ _03407_ _03408_ _03410_ _04005_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10874_ _03926_ _03929_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12613_ _05688_ _05701_ _05699_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12544_ _05755_ _05760_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12475_ _05359_ _05684_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11426_ _04042_ _04043_ _04045_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__or3_1
X_11357_ _00850_ _00821_ _01410_ _01397_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nand4_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10308_ _02581_ _02655_ _02654_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _03900_ _03896_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__and2b_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _03230_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07450_ net252 net10 VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07381_ _06145_ _06249_ _00283_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__and3_1
X_09120_ net254 net11 net13 _03820_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09051_ _01937_ _01949_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08002_ _00901_ _00902_ _00468_ _00470_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap286 _01714_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_1
X_09953_ _02917_ _02918_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__nand3_4
Xmax_cap297 _00137_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
X_08904_ _01227_ _01239_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__and2_1
X_09884_ _02840_ _02841_ _02842_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a21oi_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _01178_ _01199_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__a21bo_2
X_08766_ net223 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07717_ _00616_ _00618_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__xnor2_1
X_08697_ _01012_ _01014_ _01016_ _01001_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a22o_1
X_07648_ _02789_ _03106_ _00549_ _00550_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__nand4_2
XFILLER_0_95_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07579_ _03337_ _00058_ _00481_ net182 VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__a22o_1
X_09318_ _05115_ _01567_ _02221_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a22o_1
X_10590_ _03602_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09249_ _02146_ _02147_ _02141_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ _05449_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nand2_2
X_11211_ _03750_ _03762_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__and2b_1
X_12191_ _01563_ _03499_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__nand2_1
X_11142_ _03666_ _03669_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nor2_1
Xinput110 data_in[199] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
X_11073_ _03578_ _03582_ _03581_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__a21bo_1
Xinput143 data_in[228] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xinput121 data_in[208] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
Xinput154 data_in[238] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xinput132 data_in[218] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
X_10024_ _02981_ _02996_ _02997_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__and3_1
Xinput165 data_in[248] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
Xinput187 data_in[37] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_2
Xinput176 data_in[27] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
Xinput198 data_in[47] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11975_ net261 _05136_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10926_ _03397_ _03399_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10857_ _03910_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _03815_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__xor2_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12527_ _05735_ _05743_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or2_1
X_12458_ _02239_ _02904_ _05667_ _05413_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _04507_ _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__xor2_2
XFILLER_0_78_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12389_ _05590_ _04897_ _05591_ _01987_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06950_ net27 VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__clkbuf_4
X_06881_ _06167_ _06168_ _06194_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _03546_ _00956_ _01520_ _02635_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08551_ _01448_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08482_ _03853_ _00830_ _01380_ _01381_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__nand4_2
X_07502_ _00403_ _00404_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07433_ _00287_ _00288_ _00334_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09103_ _01981_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__xor2_2
X_07364_ _06142_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07295_ _00197_ _06281_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09034_ _01333_ _01335_ _01932_ _01933_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09936_ _02898_ _02900_ _02892_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__a21oi_1
X_09867_ _02819_ _02820_ _02824_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__o211a_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _02093_ _02095_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__or2_1
X_08818_ _01134_ _01718_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__xnor2_1
X_08749_ _01071_ _01089_ _01090_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__or3_4
XFILLER_0_95_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _04445_ _04449_ _04900_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__and3_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _02500_ _03166_ _03168_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__a21o_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _04824_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__nor2_1
X_10642_ _03051_ _03052_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ _03571_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__xor2_4
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer9 _00119_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12312_ _05497_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12243_ _05078_ _05090_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12174_ _01520_ _01484_ _02164_ _02132_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__nand4_4
X_11125_ _04165_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__xnor2_4
X_11056_ _03555_ _03560_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and2_1
X_10007_ _02318_ _02320_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11958_ _04762_ _05119_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10909_ _03966_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__or2_1
X_11889_ _00507_ _04123_ _04640_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07080_ _06392_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07982_ _00881_ _00882_ _00880_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09721_ _02663_ _02664_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__and2b_1
X_06933_ _06244_ _06245_ _06246_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__o21a_1
X_09652_ net142 net153 net154 _06177_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__a22o_1
X_06864_ _02394_ _06178_ _04150_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__nand3b_1
X_06795_ _06077_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__clkbuf_4
X_09583_ _02495_ _02511_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand3_1
X_08603_ _01501_ _01502_ _01498_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__a21o_1
X_08534_ net52 _00397_ net64 net51 VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08465_ net235 net208 net250 _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__and4_1
XFILLER_0_58_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07416_ _00315_ _00316_ _00317_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__a21o_1
X_08396_ _06178_ _01293_ _01295_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07347_ net28 VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__buf_2
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ _01915_ _01916_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07278_ _06148_ _06251_ _00180_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__nor3_1
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09919_ _02880_ _02881_ _02183_ _02853_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__o211ai_1
X_12861_ _06101_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__clkbuf_1
X_11812_ _04515_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__xnor2_2
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12792_ _05964_ _05955_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__and2b_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11743_ _04880_ _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11674_ _04354_ _04361_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__nor2_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10625_ _03569_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10556_ net230 net222 VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10487_ _02920_ _02923_ _03504_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12226_ _05412_ _05413_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__or2_1
X_12157_ _05325_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__xnor2_1
X_11108_ _03022_ _03639_ _04186_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12088_ _05260_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__nand2_1
X_11039_ _04109_ _04110_ _04101_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06580_ net51 VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08250_ _00615_ _00618_ _00614_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__o21ba_1
X_08181_ _00548_ _00552_ _00551_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__a21bo_1
X_07201_ _00103_ _00104_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07132_ _00034_ _00035_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07063_ _06374_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput266 net266 VGND VGND VPWR VPWR data_out[17] sky130_fd_sc_hd__clkbuf_4
Xoutput277 net277 VGND VGND VPWR VPWR data_out[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07965_ _00864_ _00865_ _00818_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__o21a_1
X_09704_ _02643_ _02644_ _02611_ _01932_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__o211ai_1
X_06916_ _02328_ _06227_ _06228_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__a21oi_1
X_09635_ _02544_ _02570_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__xor2_4
X_07896_ net292 _00737_ _00795_ _00796_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06847_ _04358_ _04391_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__nand2_1
X_06778_ net252 net254 _03787_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__and3b_1
X_09566_ _02485_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__xnor2_1
X_08517_ _01405_ _01416_ _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09497_ _01780_ _01782_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08448_ _00790_ net295 _01347_ _01348_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10410_ _03388_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08379_ _00692_ _00732_ _00690_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11390_ _03997_ _04008_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10341_ _03342_ _03344_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10272_ _03266_ _03267_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nand3_1
X_12011_ _05175_ _05173_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__and2b_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12844_ _06084_ _06082_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__or2_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12775_ _06005_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__xnor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _01365_ _02626_ _01986_ _00757_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a22o_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11657_ _04771_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__xnor2_1
X_10608_ _03633_ _03635_ _03637_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11588_ _04224_ _04226_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10539_ _02929_ _02937_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12209_ _05390_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__xnor2_1
X_07750_ _00252_ _00641_ _00650_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__or3_1
X_06701_ _04851_ _05049_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__xor2_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07681_ _00581_ _00582_ _00419_ _00141_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__a211oi_4
X_09420_ _02332_ _02333_ _02327_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06632_ net122 VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__buf_2
X_09351_ _02201_ _01626_ _02257_ _02258_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06563_ net114 VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08302_ _06142_ _06261_ _06264_ _00239_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__nand4_2
X_09282_ _02160_ _02161_ _02181_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__a211o_1
X_06494_ net245 VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08233_ _01132_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08164_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08095_ _00994_ _00995_ _00986_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__o21ai_1
X_07115_ _06421_ _06422_ _06428_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07046_ _06357_ _06358_ _06342_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ _01801_ _01802_ _01894_ _01895_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a22o_2
X_07948_ net3 VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__buf_4
X_07879_ _00772_ _00773_ _00779_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o21ai_1
X_10890_ _00357_ net3 net11 net13 VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__nand4_2
X_09618_ _06283_ net126 _00201_ net127 VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__nand4_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09549_ _02474_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _05773_ _05777_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__or2_1
X_11511_ _04628_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12491_ _05681_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__xor2_2
X_11442_ _04550_ _04551_ _04552_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11373_ _04476_ _04477_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10324_ _06384_ net250 _01987_ net237 VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10255_ _02744_ _02747_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__or2_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _06284_ net101 _03173_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_100_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12827_ net267 _06068_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12758_ _02174_ _05994_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11709_ _04455_ _04489_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12689_ _05919_ _05869_ _05858_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08920_ net27 net19 net20 net26 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08851_ _01749_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__or2_2
X_07802_ _04292_ _00238_ _00703_ _02251_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__a22o_1
X_08782_ _01680_ _01681_ _01649_ _01650_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__o211ai_4
X_07733_ _00337_ _00339_ _00633_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__nor3_1
X_07664_ _00563_ _00564_ _00566_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__and3_2
XFILLER_0_79_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09403_ _02312_ _02313_ _02314_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nand3_1
X_06615_ _02459_ _04106_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07595_ _00497_ _00055_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09334_ net191 net192 net188 _02239_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__nand4_2
XFILLER_0_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06546_ _03337_ _02712_ _03348_ _02723_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09265_ net78 net113 net181 VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__and3_1
X_06477_ _02558_ _02591_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09196_ _02093_ _02094_ _02060_ _02061_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08216_ net287 _01116_ _00587_ _00589_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08147_ _00536_ _00537_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08078_ _05191_ _00062_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07029_ net53 VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10040_ _01666_ _03014_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_98_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11991_ _04769_ _04789_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10942_ _02773_ _03409_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10873_ _03927_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12612_ _05833_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12543_ _05756_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12474_ _05359_ _05684_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nand2_1
X_11425_ _04034_ _04033_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11356_ _00821_ _01410_ _01397_ _00850_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__a22o_1
X_10307_ _03250_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _03936_ _03979_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21boi_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _06151_ _01872_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10169_ _03135_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__xor2_4
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ _00281_ _00282_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09050_ _01947_ _01948_ _01942_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08001_ _00468_ _00470_ _00901_ _00902_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09952_ _02217_ _02226_ _02225_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap287 _01115_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_1
Xmax_cap298 _00866_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_2
X_08903_ _01245_ _01278_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09883_ _02840_ _02841_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__and3_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _01200_ _01176_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__or2b_1
X_08765_ net212 VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07716_ net157 _00617_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08696_ _01552_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__xor2_1
X_07647_ net201 VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__buf_6
XFILLER_0_95_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07578_ _00480_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__buf_2
X_06529_ _03150_ _03161_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nor2_2
X_09317_ _00047_ _00989_ net186 _00480_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09248_ _02141_ _02146_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09179_ _02063_ _02077_ _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11210_ _03794_ _03810_ _03807_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__a21o_1
X_12190_ _01524_ _02215_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11141_ _03915_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 data_in[19] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
Xinput100 data_in[18] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
X_11072_ _04146_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__nor2_1
Xinput144 data_in[229] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xinput122 data_in[209] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
Xinput133 data_in[219] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
X_10023_ _02994_ _02995_ _02986_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__o21ai_1
Xinput166 data_in[249] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_4
Xinput155 data_in[239] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xinput177 data_in[28] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_4
Xinput199 data_in[48] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xinput188 data_in[38] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_4
XFILLER_0_98_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11974_ net261 _05136_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10925_ _03434_ _03448_ _03446_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10856_ _03906_ _03909_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__and2_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10787_ _03829_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12526_ _05737_ _05738_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12457_ _01584_ _01562_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11408_ _04508_ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12388_ _01385_ _02694_ _01367_ _02695_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11339_ _03943_ _03958_ _03957_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06880_ _06167_ _06168_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__and3_1
X_08550_ _00879_ _01449_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__a21bo_1
X_08481_ _03853_ _00830_ _01380_ _01381_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07501_ _00402_ _00401_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__and2b_1
X_07432_ _00287_ _00288_ _00334_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09102_ _02000_ _02001_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07363_ _06260_ _06269_ _06270_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__or3_1
X_07294_ _06273_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09033_ _01930_ _01931_ _01911_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09935_ _02892_ _02898_ _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09866_ net104 _02132_ _02821_ _02823_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__nand4_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _01716_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__xnor2_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _02687_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__xor2_4
X_08748_ _01089_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__inv_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08679_ _01578_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__or2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _06130_ _02464_ _03148_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a31oi_2
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _04822_ _04823_ _04816_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10641_ _03125_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10572_ _03572_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__xor2_4
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12311_ _05504_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12242_ _05041_ _05050_ _05047_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__o21a_2
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12173_ _01484_ _02164_ _02132_ _01520_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11124_ _04202_ _04204_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__xnor2_4
X_11055_ _04126_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__xnor2_2
X_10006_ _02948_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11957_ _05117_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__and2b_1
X_10908_ _06343_ _03967_ _03964_ _03965_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_98_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11888_ _04147_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10839_ _03889_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12509_ _05721_ _05722_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07981_ _00880_ _00881_ _00882_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__nand3_1
X_09720_ _02661_ _02662_ _02105_ _02107_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06932_ _04227_ _06130_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06863_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__buf_2
X_09651_ _06177_ net142 _01288_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__and3_1
X_06794_ net202 VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__clkbuf_4
X_09582_ _02496_ _02497_ _02510_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__nand3_1
X_08602_ _01498_ _01501_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__nand3_1
X_08533_ net65 VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08464_ net206 VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_4
X_07415_ _00315_ _00316_ _00317_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__nand3_1
X_08395_ _06171_ _06311_ _06319_ _00291_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__nand4_4
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07346_ net15 net28 _00247_ _00248_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09016_ _01912_ _01913_ _01914_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07277_ _00178_ _00179_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09918_ _02183_ _02853_ _02880_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__a211o_1
X_09849_ _02801_ _02804_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__nand3_1
X_12860_ _02174_ _06098_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__and3_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04955_ _04956_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _06029_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nand2_1
X_11742_ _04382_ _04425_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a21oi_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11673_ _03817_ _03826_ _04339_ _04341_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__a22o_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10624_ _03653_ _03655_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10555_ _04741_ _00086_ net224 _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nand4_2
XFILLER_0_106_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10486_ _03501_ _03503_ _03487_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__a21oi_2
X_12225_ _01617_ _01603_ _03580_ _04123_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _05335_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__nor2_1
X_11107_ _04182_ _04184_ _04185_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12087_ _05241_ _04907_ _05259_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__or3_1
X_11038_ _04101_ _04109_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__nand3_2
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08180_ _01079_ _01080_ _01078_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__a21o_1
X_07200_ _04884_ _00102_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07131_ _06436_ _00033_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07062_ _03798_ _05914_ _03831_ _06375_ _02470_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput267 net267 VGND VGND VPWR VPWR data_out[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput278 net278 VGND VGND VPWR VPWR data_out[2] sky130_fd_sc_hd__clkbuf_4
X_07964_ _00818_ _00864_ _00865_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09703_ _02611_ _01932_ _02643_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06915_ _02328_ _06227_ _06228_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__and3_1
X_07895_ net292 _00737_ _00795_ _00796_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__or4bb_1
X_09634_ _02559_ _02568_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06846_ _06158_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06777_ _02481_ _05882_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__nand2_1
X_09565_ _02491_ _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__nor2_1
X_08516_ _01414_ _01415_ _00876_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_78_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09496_ _01799_ _01801_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08447_ _01345_ _01346_ _01284_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08378_ _01245_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07329_ _04292_ _04424_ _06159_ _06134_ _06257_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10340_ _05969_ _02695_ _03343_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__and3_2
XFILLER_0_104_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10271_ _02596_ _02598_ _02597_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12010_ _05173_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__and2b_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _06084_ _06082_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__nand2_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12774_ _06006_ _06011_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__xnor2_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _04861_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__or2_2
XFILLER_0_96_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11656_ _04773_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10607_ _03633_ _03635_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11587_ _04293_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10538_ _03553_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12208_ _05391_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__xnor2_1
X_10469_ _02854_ _02878_ _02879_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nand3_1
X_12139_ _05294_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__xor2_2
X_06700_ _05016_ _05038_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__xnor2_2
X_07680_ _00419_ _00141_ _00581_ _00582_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__o211a_1
X_06631_ net86 VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09350_ _02233_ _02234_ _02255_ _02256_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06562_ _03524_ net113 net114 VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08301_ _06261_ _06264_ net19 _06142_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09281_ _02179_ _02180_ _02162_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08232_ _00603_ _00600_ _01126_ _00599_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06493_ _02756_ _02767_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08163_ _01049_ _01050_ _01064_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08094_ _00986_ _00994_ _00995_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__or3_1
X_07114_ _06426_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__xnor2_1
X_07045_ _06342_ _06357_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__and3_2
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ _01801_ _01802_ _01894_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__nand4_4
X_07947_ _00845_ _00846_ _00847_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07878_ _00772_ _00773_ _00779_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__or3_2
X_09617_ net126 net135 net127 net133 VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__a22o_1
X_06829_ _06142_ _06143_ _04479_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09548_ _01787_ _01789_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11510_ _04625_ _04627_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09479_ _01132_ _01133_ _01718_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12490_ _05682_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11441_ _04550_ _04551_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11372_ _00387_ _03967_ _02731_ _00822_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__a22oi_2
X_10323_ _06384_ net249 _02689_ _02688_ _01385_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10254_ _02650_ _02652_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__or2_1
X_10185_ net90 net98 net91 net99 VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12826_ net267 _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _05987_ _05993_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11708_ _04486_ _04488_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12688_ _05359_ _05684_ _05867_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11639_ _04335_ _04345_ _04343_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08850_ _01747_ _01748_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__and2_1
X_07801_ net99 VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_4
X_08781_ _01649_ _01650_ _01680_ _01681_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__a211o_4
X_07732_ _00337_ _00339_ _00633_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o21a_1
X_07663_ _02811_ _00107_ _00122_ _00565_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a31o_1
X_06614_ net209 VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__buf_2
X_09402_ _02312_ _02313_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09333_ net189 VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__clkbuf_4
X_07594_ _05126_ _05147_ _00051_ _00052_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06545_ net192 VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06476_ _02569_ _02580_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09264_ net110 VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09195_ _02060_ _02061_ _02093_ _02094_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08215_ _00587_ _00589_ net287 _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__a211o_2
XFILLER_0_132_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08146_ _00542_ _00567_ _00568_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08077_ _00977_ _00978_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__nor2_1
X_07028_ _02668_ _03612_ _05575_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold11 net275 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _01264_ _01265_ _01267_ _01268_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__o2bb2ai_1
X_11990_ _01777_ _01754_ _04749_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10941_ _03998_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__xor2_2
X_10872_ net238 _00834_ net250 net251 VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12611_ _05664_ _05675_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__o21a_2
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12542_ _05757_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__nor2_1
X_12473_ _02164_ _02132_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__and3_1
X_11424_ _04135_ _04094_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11355_ _04456_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11286_ _03978_ _03976_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__or2b_1
X_10306_ _03252_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10237_ _04314_ _01264_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__nand2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ _03136_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__xnor2_4
X_10099_ _02412_ _02449_ _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _06040_ _06042_ _06038_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08000_ net298 _00867_ _00899_ _00900_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09951_ _02915_ _02916_ _02907_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap299 _00573_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
X_08902_ _01799_ _01800_ _01770_ _01771_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap288 net322 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_1
X_09882_ _02141_ _02147_ _02146_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a21bo_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _01201_ _01281_ _01732_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__o21ba_2
X_08764_ net12 _00550_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07715_ net171 VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__buf_2
X_08695_ _01581_ _01595_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__xor2_1
X_07646_ net190 VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07577_ net195 VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_4
X_06528_ net41 _03084_ _03117_ _03139_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__a22oi_2
X_09316_ _00989_ net186 net195 net185 VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09247_ _02144_ _02145_ _01522_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06459_ _02383_ _02394_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09178_ _02070_ _02071_ _02076_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08129_ _01027_ _01028_ _01029_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11140_ _04220_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__xor2_4
Xinput101 data_in[190] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
X_11071_ _00086_ net230 net224 _03580_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__and4_1
Xinput134 data_in[21] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xinput145 data_in[22] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_4
Xinput123 data_in[20] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xinput112 data_in[1] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_4
X_10022_ _02986_ _02994_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__or3_1
Xinput178 data_in[29] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_4
Xinput167 data_in[24] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
Xinput156 data_in[23] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_2
Xinput189 data_in[39] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_2
XFILLER_0_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11973_ _05130_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__xor2_1
X_10924_ _03404_ _03417_ _03984_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10855_ _03906_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10786_ _03830_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _05138_ _05739_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__a21oi_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12456_ _05443_ _05447_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12387_ _02695_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__inv_2
X_11407_ _04513_ _04514_ _04515_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11338_ _03925_ _03932_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11269_ _04355_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07500_ _00401_ _00402_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__nor2b_1
X_08480_ _05980_ _06384_ _06383_ _00366_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__nand4_4
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07431_ _00331_ _00333_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ _06292_ _00263_ _00195_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__and3_1
X_09101_ _01998_ _01999_ _01984_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07293_ _06289_ _06288_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__or2b_1
X_09032_ _01911_ _01930_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__or3_2
XFILLER_0_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09934_ _02896_ _02897_ _02893_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__a21o_1
X_09865_ net104 net120 _02821_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a22o_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _00612_ _01122_ _01121_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__o21bai_2
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _02744_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_4
X_08747_ _01646_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__nand2_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08678_ _01575_ _01576_ _01577_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__a21oi_1
X_07629_ _03084_ _00097_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__nand2_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ _03671_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__xor2_2
XFILLER_0_91_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10571_ _03589_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12310_ _05499_ _05500_ _05503_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__and3_1
X_12241_ _05427_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_133_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _04539_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__xnor2_1
X_11123_ _03619_ _03648_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11054_ _05093_ _02239_ _04127_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__and3_1
X_10005_ _02949_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11956_ _05113_ _05116_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nand2_1
X_10907_ net66 VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__buf_2
X_11887_ _04642_ _04645_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10838_ _06304_ _01986_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10769_ _03255_ _03275_ _03274_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12508_ _05721_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12439_ _05643_ _05401_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07980_ _03743_ _05761_ _06343_ _00387_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__nand4_2
X_06931_ _02317_ _04238_ _06127_ _06243_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09650_ _01311_ _01909_ _01908_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__a21o_1
X_06862_ net141 VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__clkbuf_4
X_08601_ _05389_ _00438_ _01499_ _01500_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__nand4_2
X_06793_ _05871_ _06055_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__xor2_2
X_09581_ _02496_ _02497_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08532_ _00880_ _00881_ _00882_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__a21bo_1
X_08463_ net235 net249 _00828_ _00827_ _06383_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__a32o_1
X_07414_ net139 net152 VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08394_ net142 _06319_ _00291_ _06171_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__a22o_1
X_07345_ net16 _06138_ _06142_ _06264_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07276_ _06229_ _00177_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09015_ _01912_ _01913_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09917_ _02878_ _02879_ _02854_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21oi_1
X_09848_ _06424_ _00937_ _02802_ _02803_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__nand4_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _00357_ _00822_ _02726_ _02727_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand4_4
X_11810_ _01487_ _02064_ _04953_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__a21o_1
X_12790_ _06026_ _06028_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nand2_1
X_11741_ _04384_ _04423_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__nor2_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _04803_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10623_ _02979_ _03036_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10554_ net225 VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10485_ _03487_ _03501_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__and3_1
X_12224_ _01603_ _03580_ _04123_ _01617_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__a22oi_1
X_12155_ _05326_ _04984_ _05333_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__and3_1
X_11106_ _04182_ _04184_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21o_1
X_12086_ _05241_ _04907_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__o21ai_1
X_11037_ _04105_ _04107_ _04108_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11939_ _05096_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07130_ _06436_ _00033_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07061_ net255 VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput268 net268 VGND VGND VPWR VPWR data_out[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput279 net279 VGND VGND VPWR VPWR data_out[3] sky130_fd_sc_hd__clkbuf_4
X_07963_ _00862_ _00863_ _00819_ _00820_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__o211a_1
X_09702_ _02641_ _02642_ _02621_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__o21a_1
X_07894_ net295 _00793_ _00794_ _00329_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06914_ _02328_ _06130_ _06128_ _04259_ _06127_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__a32o_1
X_09633_ _02566_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__xnor2_1
X_06845_ _02240_ _06159_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09564_ _02489_ _02490_ _02486_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__a21oi_1
X_06776_ net8 VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__clkbuf_4
X_08515_ _01414_ _01415_ _00876_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__or3b_1
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09495_ _01751_ _01752_ _01757_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__o21ai_4
X_08446_ _01284_ _01345_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__or3_1
X_08377_ _01276_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07328_ _00229_ _00230_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__nor2_1
Xwire307 _00069_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__buf_1
XFILLER_0_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07259_ _00160_ _00161_ net279 VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__a21o_1
X_10270_ _03263_ _03264_ _03265_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12842_ net270 VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__inv_2
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _06009_ _06010_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__nor2_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04852_ _04853_ _04860_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__nor3_1
XFILLER_0_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _04310_ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10606_ net12 net234 _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ _04709_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10537_ _03555_ _03560_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10468_ _03483_ _03484_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or2_2
X_12207_ _01667_ _03006_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10399_ net70 net71 net83 net84 VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__nand4_2
X_12138_ _05315_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__nand2_1
X_12069_ _04894_ _04903_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nor2_1
X_06630_ _04249_ _04270_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06561_ net104 VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09280_ _02162_ _02179_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__and3_1
X_06492_ _02712_ _02723_ _02734_ _02745_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__and4_1
X_08300_ _01176_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08231_ _01125_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08162_ _01054_ _01063_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08093_ _00992_ _00993_ _00987_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a21oi_1
X_07113_ _03579_ _05520_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__nand2_1
X_07044_ _06353_ _06356_ _05838_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08995_ _01892_ _01893_ _01276_ _01803_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__a211o_1
X_07946_ _00845_ _00846_ _00847_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__a21o_1
X_07877_ _00776_ _00777_ _00778_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__or3_1
X_09616_ net124 _00665_ _01861_ _01862_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__and4_1
X_06828_ _02207_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__nand2_1
X_09547_ _02472_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__or2_2
X_06759_ _05356_ _05367_ _05685_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__or3_2
XFILLER_0_93_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09478_ _01716_ _01717_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__and2b_1
X_08429_ _01321_ _01328_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nand3_1
XFILLER_0_53_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11440_ _04038_ _04041_ _04039_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a21bo_1
X_11371_ _00387_ _00822_ _03967_ _02731_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__and4_1
X_10322_ _02693_ _02702_ _02700_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10253_ _03158_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__xnor2_4
X_10184_ _00238_ net91 net99 net90 VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12825_ _06050_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__xnor2_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _05987_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11707_ _04388_ _04421_ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a21o_2
XFILLER_0_72_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _05837_ _05846_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11638_ _04766_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11569_ _04165_ _04206_ _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08780_ _01678_ _01679_ _01659_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__a21oi_2
X_07800_ _00700_ _00701_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__nand2_1
X_07731_ net303 _00632_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07662_ _00108_ _00119_ _00120_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__and3_1
X_09401_ net44 net37 VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__and2_1
X_07593_ _00494_ _00495_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__xnor2_2
X_06613_ _04062_ _04073_ _02976_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09332_ net192 net188 net189 net191 VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a22o_1
X_06544_ net183 VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06475_ net50 VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__clkbuf_4
X_09263_ _03546_ net109 VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09194_ net305 _02092_ _02062_ _01482_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08214_ net289 _00802_ _01113_ _01114_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__o22a_1
X_08145_ _00567_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08076_ net174 net175 net111 net123 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__and4_1
X_07027_ _06122_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__inv_2
Xhold12 net276 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _01875_ _01876_ _01290_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__a21o_1
X_07929_ _02503_ _00830_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ _04000_ _04001_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__or3_2
XFILLER_0_97_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10871_ _00834_ _01367_ _01987_ _06384_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a22oi_1
X_12610_ _05660_ _05662_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12541_ _05502_ _05534_ _05537_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__nor3_1
XFILLER_0_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12472_ _01520_ _01484_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11423_ _04097_ _04134_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11354_ _00366_ _00830_ _02694_ _02695_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11285_ _03857_ _03902_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__a21bo_1
X_10305_ _03253_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__xnor2_2
X_10236_ _04128_ net155 _02589_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__a31o_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10167_ _03138_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__xnor2_2
X_10098_ _02450_ _02411_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__or2b_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12808_ _06047_ _06048_ _06049_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__o21ba_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _05973_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09950_ _02907_ _02915_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08901_ _01770_ _01771_ _01799_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__o211ai_4
Xmax_cap289 _00801_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_1
XFILLER_0_57_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09881_ _02838_ _02839_ _02830_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21o_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _01279_ _01280_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__and2b_1
X_08763_ _01660_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__xnor2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07714_ _00614_ _00615_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__nor2_1
X_08694_ _01593_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__xnor2_1
X_07645_ net179 net12 VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07576_ net123 VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06527_ net41 _03084_ _03117_ _03139_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__and4_2
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09315_ net183 _01567_ _01568_ _01569_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__and4_1
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06458_ net139 VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__clkbuf_4
X_09246_ _01522_ _02144_ _02145_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09177_ _02070_ _02071_ _02076_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a21o_1
X_08128_ _01027_ _01028_ _01029_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08059_ _00959_ _00960_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11070_ _00516_ _01617_ _03580_ _00086_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__a22oi_1
Xinput102 data_in[191] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_2
X_10021_ _02991_ _02992_ _02993_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__a21oi_1
Xinput135 data_in[220] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_4
Xinput113 data_in[200] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
Xinput124 data_in[210] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
Xinput168 data_in[250] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_2
Xinput157 data_in[240] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_2
Xinput146 data_in[230] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xinput179 data_in[2] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11972_ _03065_ _04237_ _05131_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__a31o_4
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10923_ _03412_ _03416_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__or2_1
X_10854_ _03250_ _03307_ _03907_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ _06151_ _01872_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12524_ net262 _05482_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__nor2_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12455_ _05445_ _05446_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__or2b_1
X_11406_ _03999_ _04511_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12386_ _05350_ _05387_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a21o_1
X_11337_ _03933_ _03924_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11268_ _04361_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__and2_1
X_10219_ _06274_ _01250_ _03210_ _06152_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__a22oi_1
X_11199_ _04285_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nor2_2
XFILLER_0_89_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07430_ _00332_ _06331_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07361_ _06292_ _00195_ _00263_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09100_ _01984_ _01998_ _01999_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__and3_2
XFILLER_0_57_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09031_ _01927_ _01928_ _01929_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07292_ _04358_ _06161_ _06288_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09933_ _02893_ _02896_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09864_ net105 net106 net118 net119 VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nand4_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _01714_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__or2b_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _02033_ _02051_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__a21oi_2
X_08746_ _01644_ _01645_ _01628_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__o21ai_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08677_ _01575_ _01576_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__and3_1
X_07628_ _02822_ _00530_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__nand2_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07559_ _00067_ net307 _00460_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ _03594_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__xor2_4
XFILLER_0_91_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09229_ net75 _02127_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12240_ _05074_ _05095_ _05428_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _04990_ _04991_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_102_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11122_ _03644_ _03647_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11053_ _03556_ _03558_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__or2b_1
X_10004_ _02966_ _02975_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11955_ _05113_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10906_ _06343_ net66 _03964_ _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__and4_2
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11886_ _04612_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__xor2_4
XFILLER_0_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10837_ _06173_ _01365_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10768_ _03225_ _03812_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12507_ _05178_ _05471_ _05470_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12438_ _05644_ _05057_ _05645_ _03006_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__o211a_1
X_10699_ _03700_ _03737_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__xor2_2
XFILLER_0_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12369_ _01986_ _03859_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06930_ _04238_ _06127_ _06243_ _02317_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06861_ _06174_ _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nor2_1
X_08600_ _05389_ _00438_ _01499_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a22o_1
X_06792_ _05958_ _06045_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09580_ _02501_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__xor2_1
X_08531_ _00887_ _00889_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__nand2_1
X_08462_ _00832_ _01361_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07413_ net141 net150 net151 net140 VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08393_ _04128_ _01293_ _00742_ _00743_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07344_ net17 net26 net27 net16 VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07275_ _06229_ _00177_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09014_ _03941_ net215 VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09916_ _02854_ _02878_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__and3_1
X_09847_ _06424_ _00937_ _02802_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__a22o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _00357_ _00822_ _02726_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a22o_1
X_08729_ _02822_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04844_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__xnor2_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11671_ _04792_ _04793_ _04802_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10622_ _03035_ _03033_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10553_ net229 net224 net225 net228 VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10484_ _03498_ _03500_ _03488_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12223_ _05064_ _05065_ _05069_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__a21bo_1
X_12154_ _05326_ _04984_ _05333_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__a21oi_1
X_11105_ _01666_ net45 VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__and2_1
X_12085_ _05247_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__xor2_2
X_11036_ _04105_ _04107_ _04108_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__nand3_2
XFILLER_0_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11938_ _04657_ _04691_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11869_ _05001_ _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07060_ _05914_ _03787_ _06373_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput258 net258 VGND VGND VPWR VPWR data_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput269 net269 VGND VGND VPWR VPWR data_out[1] sky130_fd_sc_hd__clkbuf_4
X_09701_ _02621_ _02641_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__nor3_1
X_07962_ _00819_ _00820_ _00862_ _00863_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__a211oi_2
X_07893_ _00329_ _00792_ _00793_ _00794_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__or4_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06913_ net169 VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__clkbuf_4
X_09632_ _01878_ _01879_ _01877_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__a21boi_1
X_06844_ net87 VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__clkbuf_4
X_09563_ _02486_ _02489_ _02490_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__and3_1
X_08514_ _01408_ _01409_ _01411_ _01413_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__a22oi_2
X_06775_ _03842_ _03908_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09494_ _01894_ _01896_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__nand2_4
X_08445_ _01343_ _01344_ _00864_ _00866_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08376_ _01246_ _00688_ _01275_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07327_ net86 _06253_ _00227_ _00228_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07258_ net279 _00160_ _00161_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__nand3_1
X_07189_ _04818_ _00092_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12841_ _06083_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _05923_ _06007_ _06008_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__and3_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _04852_ _04853_ _04860_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _04783_ _04784_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__or2_1
X_10605_ _03106_ net223 VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11585_ _03915_ _04223_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10536_ _03556_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10467_ _03481_ _03482_ _03450_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a21oi_1
X_12206_ _01666_ _01652_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10398_ _06424_ _01443_ _02064_ _05498_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__a22o_1
X_12137_ _05314_ _05295_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _04864_ _04875_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__o21ba_2
X_11019_ _04087_ _04088_ _04024_ _04025_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06560_ _02899_ _03502_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06491_ _02712_ _02723_ _02734_ _02745_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08230_ _00166_ _01131_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__nor2_1
X_08161_ _01061_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__nor2_1
X_07112_ _06423_ _06425_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__or2b_1
X_08092_ _00987_ _00992_ _00993_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07043_ _05838_ _06353_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__or3_2
XFILLER_0_70_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08994_ _01276_ _01803_ _01892_ _01893_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07945_ net253 net10 VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07876_ _00292_ _00775_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__nor2_2
X_09615_ net125 _06283_ _00210_ _00201_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06827_ net26 VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__clkbuf_4
X_09546_ _02471_ net31 _04435_ _02468_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__and4b_1
X_06758_ _05663_ _05674_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__or2_1
X_09477_ _02396_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__nor2_1
X_08428_ _01326_ _01327_ _01322_ _01323_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a211o_1
X_06689_ net1 net12 VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08359_ _00667_ _00669_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11370_ _03988_ _03994_ _03993_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__a21oi_2
X_10321_ _02673_ _02678_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10252_ _03245_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__nor2_2
X_10183_ _02499_ _02500_ _02509_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__nor3_1
X_12824_ _06056_ _06065_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12755_ _05988_ _05989_ _05990_ _05737_ _05992_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__a221o_1
X_11706_ _04422_ _04386_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__and2b_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _05845_ _05839_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__and2b_1
X_11637_ _04301_ _04316_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2b_1
XFILLER_0_107_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11568_ _04202_ _04204_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10519_ _03537_ _03538_ _03539_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11499_ _04615_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07730_ _00630_ _00631_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ _02811_ _00543_ _00561_ _00562_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a22o_1
X_09400_ _03194_ net43 _01068_ net39 VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nand4_1
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07592_ _02712_ _03348_ _05115_ _00049_ _00052_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a41o_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06612_ _02976_ _04062_ _04073_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nand3_2
X_09331_ _05093_ _00489_ _01586_ _01585_ _01584_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__a32o_1
X_06543_ _03304_ _03315_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06474_ net59 VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09262_ _01529_ _01531_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09193_ _02062_ _01482_ net305 _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08213_ net289 _00802_ _01113_ _01114_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__nor4_1
X_08144_ _01022_ _01045_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08075_ _05202_ _00059_ _00479_ _03392_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07026_ _06337_ _06338_ _06192_ _06242_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__o211a_1
X_08977_ _01290_ _01875_ _01876_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__nand3_1
X_07928_ net249 VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_4
X_07859_ _04106_ _06077_ _06172_ _06361_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__and4_1
X_10870_ _03336_ _03339_ _03338_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09529_ _01795_ _01797_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__and2_2
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12540_ _05534_ _05537_ _05502_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__o21a_2
XFILLER_0_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12471_ _05431_ _05451_ _05449_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_53_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11422_ _04085_ _04087_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__or2b_2
XFILLER_0_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11353_ _00830_ _02694_ _02695_ _00366_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11284_ _03903_ _03855_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2b_1
X_10304_ _03254_ _03303_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10235_ _06177_ net142 net153 net154 VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__and4_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ _03151_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10097_ _03057_ _02409_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12807_ _06047_ _06048_ _00166_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__a21o_1
X_10999_ _04065_ _04066_ _04067_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05749_ _05895_ _05894_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12669_ _05897_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08900_ _01797_ _01798_ _01772_ _01243_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__a211o_1
X_09880_ _02830_ _02838_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__nand3_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08831_ _06229_ _00177_ _00625_ _01166_ _01164_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a41o_2
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _01661_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__and2b_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _01013_ _01010_ _01011_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__o21ai_1
X_07713_ net159 _06227_ _00171_ _04227_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__a22oi_2
X_07644_ _00545_ _00546_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07575_ _00476_ _00477_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06526_ _02800_ _03128_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__nand2_4
XFILLER_0_118_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09314_ net184 _00049_ _00058_ _00481_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__and4_1
X_06457_ net148 VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__clkbuf_4
X_09245_ _06437_ net117 _02142_ _02143_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09176_ _02074_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__xor2_2
XFILLER_0_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ net217 _00516_ _00519_ _00518_ _04741_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__a32o_1
X_08058_ _00954_ _00955_ _00957_ _00958_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a22o_1
X_07009_ _06181_ _06321_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nor3_2
XFILLER_0_12_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10020_ _02991_ _02992_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__and3_1
Xinput136 data_in[221] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xinput103 data_in[192] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xinput125 data_in[211] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_4
Xinput114 data_in[201] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xinput169 data_in[251] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
Xinput147 data_in[231] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xinput158 data_in[241] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_2
X_11971_ _04250_ _05132_ _05131_ _04240_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__a221o_1
X_10922_ _03450_ _03482_ _03481_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10853_ _03252_ _03306_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10784_ _03230_ _03231_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12523_ net262 _05482_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12454_ _05660_ _05662_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11405_ _04509_ _04510_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12385_ _05386_ _05352_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11336_ _04023_ _04090_ _04089_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11267_ _04359_ _04360_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__or2_1
X_10218_ net138 VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__clkbuf_4
X_11198_ _04266_ _04267_ _04284_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__and3_1
X_10149_ _02478_ _02461_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07360_ _00224_ _00262_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09030_ _01927_ _01928_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07291_ _06301_ _06335_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09932_ _02894_ _02895_ net176 _00985_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_110_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09863_ net106 net118 net119 net105 VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _02050_ _02049_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__and2b_1
X_08814_ _01712_ _01713_ _01136_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__o21ai_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _01628_ _01644_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__or3_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _00986_ _00995_ _00994_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__o21bai_1
X_07627_ net46 VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_4
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ net307 _00460_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06509_ _02690_ _02701_ _02932_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07489_ _00388_ _00389_ _00390_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09228_ net77 net74 net75 net76 VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__a22o_1
X_09159_ _01432_ _01457_ _02058_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _05026_ _05052_ _05351_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11121_ _04181_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11052_ _04122_ _04125_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__xnor2_2
X_10003_ _02973_ _02974_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11954_ _04434_ _04708_ _05114_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__a21oi_2
X_10905_ _06368_ _00822_ _01410_ _02731_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__nand4_2
X_11885_ _05037_ _05039_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__nand2_2
XFILLER_0_129_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10836_ _03887_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10767_ _03228_ _03233_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10698_ _03702_ _03736_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__xnor2_4
X_12506_ _05516_ _05720_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12437_ _01666_ _01667_ _01652_ _03019_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12368_ _05251_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__xnor2_4
X_11319_ _03883_ _03895_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a21o_1
X_12299_ _05179_ _05271_ _05492_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06860_ _03941_ _02459_ _04106_ _06173_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06791_ _03897_ _06034_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08530_ _00936_ _00948_ _00935_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__a21bo_1
X_08461_ _00371_ _00372_ _00836_ _00837_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07412_ net140 _06177_ net150 net151 VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08392_ net152 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07343_ _00245_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__inv_2
X_07274_ _00175_ _00176_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _06086_ _06361_ net213 _00757_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__nand4_1
XFILLER_0_103_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09915_ _02875_ _02876_ _02231_ net304 VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09846_ _06410_ _00431_ _00421_ _01487_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__nand4_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _05882_ _06368_ _00850_ net4 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__nand4_4
X_06989_ _02448_ _06086_ _06066_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__and3_1
X_08728_ net48 VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _00978_ _01553_ _01558_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__nor3_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _04792_ _04793_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10621_ _03600_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10552_ _03575_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12222_ _05084_ _05089_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nor2_1
X_10483_ _03488_ _03498_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__nand3_2
XFILLER_0_32_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12153_ _05330_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11104_ _00109_ _00544_ _01667_ _03019_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__nand4_1
XFILLER_0_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12084_ _05255_ _05256_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__nand2_1
X_11035_ _03537_ _03539_ _03538_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11937_ _04687_ _04690_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11868_ _05019_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nor2_1
X_10819_ _03263_ _03265_ _03264_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11799_ _04044_ _04045_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput259 net259 VGND VGND VPWR VPWR data_out[10] sky130_fd_sc_hd__clkbuf_4
X_07961_ _00842_ _00843_ _00861_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09700_ _02638_ _02639_ _02640_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06912_ _04523_ _06164_ _06166_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a21o_1
X_07892_ _00332_ _00330_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__nor2_1
X_09631_ _02560_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__xor2_1
X_06843_ _04347_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06774_ _05838_ _05849_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nand2_1
X_09562_ _00239_ _00250_ _02487_ _02488_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__nand4_2
X_08513_ _01408_ _01409_ _01411_ _01413_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09493_ _01735_ _01756_ _01757_ _01759_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__a32o_2
XFILLER_0_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08444_ _00864_ _00866_ _01343_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__o211a_2
XFILLER_0_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08375_ _01246_ _00688_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07326_ _04292_ _06253_ _00227_ _00228_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07257_ _00158_ _00159_ _06224_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07188_ _00090_ _00091_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09829_ _02751_ _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__xor2_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12840_ _02174_ _06081_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__and3_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12771_ _05923_ _06007_ _06008_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a21oi_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _04854_ _04859_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__xnor2_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _04781_ _04782_ _03772_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__a21oi_1
X_10604_ _03630_ _03631_ _03632_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11584_ _04220_ _04222_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10535_ net193 _02239_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10466_ _03450_ _03481_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__and3_1
X_12205_ _01652_ _03019_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10397_ _03405_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__nor2_1
X_12136_ _05295_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12067_ _04872_ _04874_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__and2b_1
X_11018_ _04024_ _04025_ _04087_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06490_ net78 VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08160_ _01058_ _01059_ _01060_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07111_ net77 _05498_ _06424_ net76 VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08091_ _00990_ _00991_ _00988_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07042_ _06354_ _06355_ _05783_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08993_ _01849_ _01850_ _01890_ _01891_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__a2bb2o_1
X_07944_ _05914_ _05882_ _06375_ _06368_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__nand4_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07875_ _04139_ _00291_ _00774_ _02383_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__a22oi_1
X_09614_ _02545_ _02546_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nor2_1
X_06826_ _06139_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09545_ _04435_ _01784_ _02469_ _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__o2bb2a_1
X_06757_ _05378_ _05652_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__and2_1
X_06688_ _02811_ _04906_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09476_ _02393_ _02395_ _01712_ net286 VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__a211oi_1
X_08427_ _01322_ _01323_ _01326_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_108_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08358_ _01257_ _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07309_ _06152_ _06151_ _00209_ _00211_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08289_ net168 _00270_ _01187_ _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__o2bb2a_1
X_10320_ _02674_ _02677_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10251_ _03159_ _03160_ _03244_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10182_ _03168_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12823_ _06057_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12754_ _05735_ _05742_ _05901_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__and3_1
X_11705_ _04839_ _04841_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__nor2_4
XFILLER_0_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12685_ _05865_ _05876_ _05874_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11636_ _04302_ _04315_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11567_ _04657_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10518_ _03537_ _03538_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11498_ _04109_ _04111_ _04614_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10449_ _03461_ _03462_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12119_ _04915_ _04914_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__or2b_1
X_07660_ _02811_ _00543_ _00561_ _00562_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__nand4_4
X_07591_ _00492_ _00493_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__or2_1
X_06611_ _03710_ _03721_ _04051_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a21o_1
X_09330_ _01606_ _01614_ _01613_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__a21o_1
X_06542_ _02877_ _03293_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09261_ _01561_ _01578_ _01579_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06473_ _02536_ _02547_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__nand2_1
X_08212_ net321 _01112_ _00803_ _00804_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09192_ _02079_ _02080_ _02090_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08143_ _00540_ _01044_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08074_ _00473_ _00475_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07025_ _06192_ _06242_ _06337_ _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_113_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08976_ _06151_ _00677_ _01873_ _01874_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nand4_1
X_07927_ _06383_ _00827_ _00828_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__a21bo_1
X_07858_ _00758_ _00759_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07789_ _00688_ _00689_ _00662_ _00221_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__a211oi_1
X_06809_ _03710_ _04062_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09528_ _02452_ _01967_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09459_ _01695_ _02110_ _02376_ _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_54_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12470_ _05380_ _05381_ _05384_ _05680_ _05368_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a32o_1
X_11421_ _04437_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__xor2_4
XFILLER_0_62_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11352_ _04440_ _04454_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__xor2_2
XFILLER_0_131_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10303_ _03277_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11283_ _04377_ _04378_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__and2_2
X_10234_ _02560_ _02565_ _03226_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__a21o_1
X_10165_ _02491_ _03140_ _03149_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__nor3_1
X_10096_ _03055_ _03056_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12806_ _05984_ _05995_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nand2_1
X_10998_ net123 net180 VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _05970_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _05489_ _05725_ _05723_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11619_ _03717_ _04275_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__and2b_1
X_12599_ _05819_ _05820_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _01353_ _01355_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__and2_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _00549_ _00109_ _00544_ _04939_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08692_ _01582_ _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__xnor2_1
X_07712_ net158 net159 _06227_ _00171_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__and4_1
X_07643_ _03095_ _00109_ _00544_ _02800_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a22oi_1
X_09313_ _02214_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__xnor2_1
X_07574_ _00474_ _00475_ _00064_ _00066_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__o211a_1
X_06525_ net112 net245 net256 VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__and3_4
XFILLER_0_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09244_ _06437_ net117 _02142_ _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06456_ _02350_ _02361_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09175_ _06347_ _00387_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08126_ net218 _00516_ _01025_ _01026_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08057_ _00954_ _00955_ _00957_ _00958_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07008_ _04128_ net139 _06171_ _06319_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput115 data_in[202] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput104 data_in[193] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_4
Xinput126 data_in[212] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_2
Xinput159 data_in[242] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
Xinput148 data_in[232] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
Xinput137 data_in[222] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
X_08959_ net94 _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nand2_1
X_11970_ _04253_ _04718_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__nor2_1
X_10921_ _03393_ _03418_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10852_ _03850_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10783_ _06178_ _02592_ _03258_ _03257_ _00749_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__a32o_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12522_ _05138_ _05139_ _05483_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__and3_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12453_ _05403_ _05405_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11404_ _03999_ _04511_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__or2_1
X_12384_ _05318_ _05584_ _05585_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__a21bo_1
X_11335_ _03980_ _04016_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__a21o_2
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11266_ _04359_ _04360_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nand2_1
X_10217_ _03208_ _02607_ _02606_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11197_ _04266_ _04267_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a21oi_1
X_10148_ _02477_ _02463_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__or2b_1
X_10079_ _02391_ _02393_ _03058_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07290_ _06189_ _06333_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09931_ _02894_ _02895_ net176 _00985_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09862_ net103 net120 _02133_ _02134_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__and4_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _02722_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08813_ _01136_ _01712_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__nor3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _01642_ _01643_ _01069_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__o21ba_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _01573_ _01574_ _01566_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__a21o_1
X_07626_ _00106_ _00123_ _00124_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__nand3_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07557_ _00458_ _00459_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06508_ _02690_ _02701_ _02932_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07488_ _00388_ _00389_ _00390_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09227_ net76 net77 net74 VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__and3_1
X_06439_ _02174_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09158_ _01455_ _01456_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09089_ net236 net235 net250 net251 VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__and4_1
X_08109_ _00522_ _01009_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11120_ _04198_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__xor2_4
XFILLER_0_102_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11051_ _03574_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__nor2_1
X_10002_ _01619_ _02289_ _02288_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11953_ _04705_ _04707_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__nor2_1
X_10904_ _00822_ _01410_ _02731_ _06368_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a22o_1
X_11884_ _05029_ _05030_ _05036_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__nand3_1
X_10835_ _00343_ _02626_ _03884_ _03885_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__nand4_1
XFILLER_0_67_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10766_ _03228_ _03233_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10697_ _03703_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__xnor2_4
X_12505_ _05717_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12436_ _03019_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12367_ _02615_ _02592_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11318_ _03892_ _03894_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12298_ _05181_ _05270_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__or2b_1
X_11249_ _04339_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06790_ _06012_ _06023_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ _00836_ _00837_ _00371_ _00372_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08391_ _06178_ _06171_ _06311_ _06319_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__and4_1
X_07411_ _00290_ _00313_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07342_ _00243_ _00244_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07273_ _06245_ _06248_ _00174_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__or3_1
X_09012_ _06361_ net213 net214 _06077_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09914_ _02231_ net304 _02875_ _02876_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09845_ net72 _00421_ net73 _06410_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__a22o_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ net9 net3 net4 _05882_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__a22o_1
X_06988_ _05871_ _06055_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__nor2_1
X_08727_ _01054_ _01063_ _01061_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _00978_ _01553_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__o21a_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _00509_ _00510_ _00511_ _00081_ _04785_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__o32a_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _02657_ _03590_ _01487_ _01488_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__nand4_2
X_10620_ _03649_ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10551_ _04752_ net233 VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10482_ _05191_ _03499_ _03496_ _03497_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nand4_2
X_12221_ _05407_ _05088_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12152_ _01434_ _02765_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__and3_1
X_11103_ _00544_ _01667_ net234 _00109_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__a22o_1
X_12083_ _05248_ _05254_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__nand2_1
X_11034_ _04102_ _04103_ _04104_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11936_ _05074_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_129_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11867_ _05018_ _05002_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__and2b_1
X_10818_ _03867_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__nand2_1
X_11798_ _04508_ _04516_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__a21o_2
XFILLER_0_131_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10749_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12419_ _05624_ _02799_ _04953_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07960_ _00842_ _00843_ _00861_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__nor3_2
X_06911_ _04084_ _04622_ _06203_ _06204_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__a211o_1
X_07891_ _00790_ _00791_ _00327_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09630_ _02561_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__xor2_1
X_06842_ _06155_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06773_ _03765_ _05827_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__or2_1
X_09561_ _00239_ net28 _02487_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08512_ _00852_ _01412_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__xnor2_1
X_09492_ _01159_ _01160_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__and2_1
X_08443_ _01341_ _01342_ _01285_ _00784_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08374_ _01248_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__xor2_1
X_07325_ _04424_ net87 _06134_ net88 VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__nand4_1
XFILLER_0_45_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07256_ _06224_ _00158_ _00159_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__nand3_2
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07187_ _00085_ _00089_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09828_ _02752_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__xnor2_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _06375_ net11 net13 net254 VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a22o_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05940_ _05942_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__or2_2
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _04857_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__nand2_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _03772_ _04781_ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10603_ _03630_ _03631_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11583_ _04434_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10534_ _03348_ _01584_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10465_ _03477_ _03479_ _03451_ _02846_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__o211ai_2
X_12204_ _01072_ _03019_ _05061_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__and3_1
X_10396_ _05761_ net62 net57 net58 VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12135_ _05305_ _05313_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__xor2_1
X_12066_ _04908_ _04936_ _05237_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11017_ _04085_ _04086_ _04058_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11919_ _04682_ _04675_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12899_ clknet_1_1__leaf_clk _00023_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07110_ net71 VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08090_ _00988_ _00990_ _00991_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07041_ _05805_ _06352_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _01849_ _01850_ _01890_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__or4bb_4
X_07943_ net8 net255 net9 net254 VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__a22o_1
X_07874_ _00292_ _00775_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__and2_1
X_09613_ _04303_ net124 net137 net138 VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__and4_1
X_06825_ _06138_ _04468_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__and2_1
X_09544_ net17 net18 net29 net30 VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__and4_1
X_06756_ _05378_ _05652_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__nor2_1
X_06687_ net35 VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__clkbuf_4
X_09475_ _01712_ net286 _02393_ _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08426_ _06362_ _06304_ _01324_ _01325_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__nand4_1
XFILLER_0_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08357_ _04303_ _00665_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07308_ net130 net131 net125 _00210_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__nand4_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08288_ _02317_ _04238_ net162 _01188_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07239_ _06408_ _05696_ _00141_ _00142_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10250_ _03159_ _03160_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10181_ _02488_ _02490_ _03167_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12822_ _06061_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__xnor2_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _05735_ _05738_ _05901_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11704_ _04791_ _04838_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__and2_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12684_ _05910_ _05913_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__xnor2_1
X_11635_ _04437_ _04529_ _04528_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a21o_2
XFILLER_0_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11566_ _04687_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__xor2_4
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10517_ net186 net196 VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__and2_1
X_11497_ _04109_ _04111_ _04614_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10448_ _02830_ _02839_ _02838_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10379_ _02752_ _02782_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a21bo_1
X_12118_ _04920_ _04921_ _04932_ _04931_ _04929_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__o32a_1
X_12049_ _05216_ _05217_ _04856_ _04858_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o211ai_1
X_07590_ _00490_ _00491_ _05115_ _05093_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__and4bb_1
X_06610_ _03710_ _03721_ _04051_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06541_ _02877_ _03293_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__or2_1
X_06472_ _02448_ _02459_ _02514_ _02525_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__a22o_2
XFILLER_0_87_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09260_ _01575_ _01576_ _01577_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08211_ _00803_ _00804_ net321 _01112_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_117_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09191_ _02079_ _02080_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_62_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08142_ _01033_ _01043_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08073_ _00055_ _00496_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07024_ _06116_ _06119_ _06336_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08975_ _06151_ _00677_ _01873_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__a22o_1
X_07926_ net237 net247 net248 net236 VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__a22o_1
X_07857_ _03941_ _02459_ _00297_ _00757_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07788_ _00662_ _00221_ _00688_ _00689_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__o211a_1
X_06808_ _05729_ _05740_ _06121_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__o21ai_1
X_09527_ _01345_ _01898_ _01963_ _01964_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__o211a_1
X_06739_ _05455_ _05466_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09458_ _02374_ _02375_ _02197_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08409_ net149 _00774_ _01309_ _02383_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__a22o_1
X_09389_ _02298_ _02299_ _02266_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11420_ _04528_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11351_ _04441_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10302_ _03300_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11282_ _04319_ _04376_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10233_ _02561_ _02564_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__and2_1
X_10164_ _02491_ _03140_ _03149_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10095_ _03061_ _03065_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12805_ _06044_ _06046_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10997_ _00453_ net134 net178 net145 VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__nand4_1
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12736_ _05754_ _05764_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _05749_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11618_ _04744_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__or2_1
X_12598_ _05819_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11549_ _04174_ _04176_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ net179 _00549_ _00109_ _00544_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__and4_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08691_ _01583_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__xnor2_1
X_07711_ _06232_ _00187_ _00185_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__a21oi_2
X_07642_ _03095_ net1 _00109_ _00544_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__and4_1
X_09312_ net167 _02215_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nand2_1
X_07573_ _00064_ _00066_ _00474_ _00475_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a211oi_2
X_06524_ _03095_ _02789_ _03106_ _02800_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09243_ net115 net116 net107 net108 VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__nand4_2
XFILLER_0_16_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06455_ _02295_ _02306_ _02339_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09174_ _01444_ _02072_ _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08125_ _03227_ _00516_ _01025_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__nand4_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _02635_ _03546_ _00454_ _00956_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__nand4_2
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07007_ _06320_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput116 data_in[203] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_4
Xinput105 data_in[194] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
Xinput127 data_in[213] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
Xinput149 data_in[233] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
Xinput138 data_in[223] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
X_08958_ net93 VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_4
X_07909_ _02448_ _00810_ _00368_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__nand3_2
X_08889_ _01787_ _01784_ net15 _01785_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__and4b_1
X_10920_ _03419_ _03391_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__and2b_1
X_10851_ _03852_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__xor2_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10782_ _03818_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _03691_ _03692_ _04245_ _04723_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a41o_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _05406_ _05426_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__or2_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11403_ _04509_ _04510_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12383_ _05342_ _05344_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__or2b_1
X_11334_ _04013_ _04015_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__nor2_1
X_11265_ _03819_ _03822_ _03821_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10216_ _01947_ _01949_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__nand2_1
X_11196_ _04282_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__xor2_1
X_10147_ _02538_ _02540_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__nor2_2
X_10078_ _02409_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_12719_ _05815_ _05886_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09930_ net174 net175 net145 net156 VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09861_ net104 net105 _00910_ net119 VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__and4_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _02740_ _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__xnor2_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _01710_ _01711_ _01117_ _01137_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__o211a_1
X_08743_ _01642_ _01643_ _01069_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_84_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08674_ _01566_ _01573_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__nand3_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _00526_ _00527_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07556_ _02745_ _00453_ _00457_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06507_ _02899_ _02921_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07487_ net51 net62 VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__and2_1
X_09226_ _02113_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__xnor2_2
X_06438_ net257 VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09157_ _01459_ _01430_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09088_ _03853_ net250 _01987_ net235 VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__a22oi_1
X_08108_ _00522_ _01009_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08039_ _02668_ _00937_ _00938_ _00940_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11050_ _04752_ _04123_ _03575_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__and3_1
X_10001_ _02967_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ _04889_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__xnor2_2
X_10903_ _03394_ _03401_ _03400_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11883_ _05029_ _05030_ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a21o_1
X_10834_ _00343_ net215 _03884_ _03885_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10765_ _03794_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12504_ _05714_ _05716_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10696_ _03704_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ _05390_ _05394_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12366_ _05288_ _05293_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11317_ _04415_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12297_ _05152_ _05170_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__a21o_2
X_11248_ _03816_ _03817_ _03828_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__o31ai_2
X_11179_ _06243_ _01754_ _03728_ _03726_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a31o_2
X_08390_ _01289_ _01290_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nor2_1
X_07410_ _00311_ _00312_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07341_ _02251_ _00238_ _00240_ _00241_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ _06245_ _06248_ _00174_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o21ai_1
X_09011_ _01311_ _01910_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09913_ _02873_ _02874_ _02856_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__a21o_1
X_09844_ net79 _01487_ _02128_ _02127_ _02799_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__a32o_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _02081_ _02088_ _02087_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a21oi_2
X_06987_ _06299_ _06300_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__nor2_1
X_08726_ _01041_ _01602_ _01625_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nor3_1
XFILLER_0_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _01556_ _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__xnor2_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _00081_ _00508_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08588_ _03590_ _01487_ _01488_ _02657_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07539_ _02646_ _00438_ _00439_ _00440_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10550_ _03573_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09209_ _02107_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__nor2_2
X_10481_ net181 VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _05085_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12151_ _00872_ _01444_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__nand2_1
X_11102_ _04167_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__xnor2_4
X_12082_ _05248_ _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__or2_1
X_11033_ _04102_ _04103_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11935_ _05092_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11866_ _05002_ _05018_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__and2b_1
X_10817_ _06319_ _01293_ _01309_ _02615_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand4_2
X_11797_ _04507_ _04517_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10748_ _03778_ _03779_ _03790_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12418_ _01487_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__inv_2
X_10679_ _03098_ _03099_ _03097_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12349_ _04869_ _05242_ _05244_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__a21oi_1
X_06910_ _06216_ _06217_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__and2_1
X_07890_ _00327_ _00790_ _00791_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__nor3_1
X_06841_ _02229_ _06151_ _06153_ _06154_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06772_ _03765_ _05827_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__nand2_1
X_09560_ _06142_ _06264_ net20 _01217_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__nand4_2
XFILLER_0_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08511_ net6 _03798_ net3 net4 VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__and4_2
XFILLER_0_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09491_ _01969_ _01971_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__and2_2
X_08442_ _01285_ _00784_ _01341_ _01342_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08373_ _01249_ _01273_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07324_ net87 _06254_ net88 _04413_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07255_ _00156_ _00157_ _06211_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_121_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07186_ _00085_ _00089_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09827_ _02753_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__xnor2_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _02036_ _02039_ _02037_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__a21bo_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ net228 net220 _00086_ net221 VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__nand4_4
XFILLER_0_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09689_ _04106_ _06173_ net206 net207 VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__nand4_2
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _00774_ _02592_ _04855_ _04856_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand4_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _04306_ _04308_ _04780_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ _00550_ net45 VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11582_ _04705_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__xor2_4
XFILLER_0_64_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10533_ _01023_ _02950_ _02952_ _02953_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10464_ _03451_ _02846_ _03477_ _03479_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10395_ _06347_ _01444_ _02765_ _05761_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a22oi_1
X_12203_ _05350_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _05310_ _05311_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12065_ _04933_ _04935_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11016_ _04058_ _04085_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11918_ _04646_ _04651_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12898_ clknet_1_1__leaf_clk _00022_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11849_ _04996_ _04999_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__xor2_4
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07040_ _05805_ _06352_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08991_ _01888_ _01889_ _01851_ _01852_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__o211ai_2
X_07942_ _00363_ _00361_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__and2b_1
X_07873_ net148 net149 _00291_ _00774_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__and4_2
X_09612_ _06152_ net137 net138 _04303_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__a22oi_1
X_06824_ _04435_ _04446_ _06138_ _02196_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_92_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09543_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__inv_2
X_06755_ _05619_ _05641_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__or2_1
X_06686_ _04873_ _04884_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__nor2_2
X_09474_ _02391_ _02392_ _01727_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__a21o_1
X_08425_ _06362_ _06304_ _01324_ _01325_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__a22o_1
X_08356_ _01255_ _01256_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07307_ net126 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08287_ net163 VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__buf_2
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07238_ _00139_ _00140_ _00043_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__a21oi_1
X_07169_ _00057_ _00071_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__or2_1
X_10180_ _02488_ _02490_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__a21oi_1
X_12821_ _06009_ _06062_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12752_ net263 _05734_ _05900_ net264 VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__a22o_1
X_11703_ _04791_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__nor2_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05911_ _05847_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11634_ _04377_ _04378_ _04430_ _04429_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a31o_2
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11565_ _04181_ _04201_ _04689_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10516_ _00989_ _00480_ net187 net188 VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nand4_2
X_11496_ _04609_ _04613_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10447_ _03459_ _03460_ _03453_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10378_ _02753_ _02781_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__or2b_1
X_12117_ _05292_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand2_1
X_12048_ _04856_ _04858_ _05216_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__a211o_1
X_06540_ _03216_ _03282_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06471_ _02448_ _02459_ _02514_ _02525_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nand4_4
XFILLER_0_118_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08210_ _00905_ _00906_ _01109_ _01110_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__o22a_1
X_09190_ _02081_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08141_ _01041_ _01042_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08072_ _00499_ _00488_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07023_ _06116_ _06119_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08974_ _02218_ _04314_ _01264_ _01872_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07925_ net236 net237 net248 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__and3_1
X_07856_ _03941_ _00297_ _00757_ _02459_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__a22oi_1
X_07787_ _00663_ _00664_ _00687_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__nand3_1
X_06807_ _05729_ _05740_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__or3_2
XFILLER_0_78_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06738_ _05444_ _03535_ _02646_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__o21a_1
X_09526_ _02411_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__xnor2_2
X_09457_ _02197_ _02374_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08408_ net146 VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06669_ _02185_ _04688_ _04699_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__and3_1
X_09388_ _02266_ _02298_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08339_ _01227_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11350_ _04450_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10301_ _02621_ _02642_ _02641_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11281_ _04319_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_2
X_10232_ _03213_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__xor2_2
X_10163_ _03141_ _03148_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__xnor2_1
X_10094_ _02391_ _02393_ _03058_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12804_ net266 _06043_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10996_ net134 net178 net145 net177 VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a22o_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _05765_ _05752_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _05894_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12597_ _03580_ _04123_ _05654_ _05068_ _04154_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11617_ _04742_ _04743_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__and2_1
X_11548_ _04669_ _04670_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11479_ _04592_ _04593_ _04565_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _00170_ _00190_ _00189_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__o21ba_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08690_ _01589_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__xor2_1
X_07641_ net34 VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07572_ _00472_ _00473_ _03381_ _00062_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__and4bb_1
X_06523_ net256 VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__clkbuf_4
X_09311_ net156 VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09242_ net116 net107 net108 net115 VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06454_ _02295_ _02306_ _02339_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and3_2
XFILLER_0_133_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09173_ net61 net55 net57 net60 VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08124_ _04752_ _04741_ net220 _00086_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nand4_1
XFILLER_0_31_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08055_ net114 _00454_ _00956_ net113 VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__a22o_1
X_07006_ _04128_ _06171_ _06319_ _02394_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput106 data_in[195] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
Xinput117 data_in[204] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_4
Xinput139 data_in[224] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
Xinput128 data_in[214] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
X_08957_ _01855_ _01856_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nor2_1
X_07908_ net205 VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__clkbuf_4
X_08888_ net15 _01784_ _01786_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__o2bb2a_1
X_07839_ _06364_ _00347_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__nor2_1
X_10850_ _03855_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10781_ _03826_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _02428_ _02430_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _04243_ _04726_ _04722_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _05649_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__xor2_4
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11402_ net73 _01443_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12382_ _05346_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__inv_2
X_11333_ _04294_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__xor2_4
XFILLER_0_22_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11264_ _04356_ _04357_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nor2_1
X_10215_ _02559_ _03204_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__o21ai_2
X_11195_ _00270_ _01754_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10146_ _02457_ _02480_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a21bo_2
X_10077_ _03055_ _03056_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10979_ _04044_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__xor2_4
XFILLER_0_84_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12718_ _05883_ _05885_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12649_ _05865_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09860_ _02816_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _02034_ _02048_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__a21oi_4
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _01117_ _01137_ _01710_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__a211oi_4
X_08742_ _01640_ _01641_ _01634_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__a21oi_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _01570_ _01571_ _01572_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__a21o_1
X_07624_ _00506_ _00090_ _00525_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__nor3_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07555_ _02745_ _00453_ _00457_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07486_ _03743_ _05750_ _05761_ _06343_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__nand4_1
XFILLER_0_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06506_ _02778_ _02910_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09225_ _02123_ _02124_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09156_ _01458_ _01431_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09087_ net251 VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08107_ _01007_ _01008_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08038_ _00939_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10000_ _02968_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__xnor2_2
X_09989_ _02957_ _02958_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11951_ _05109_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__xor2_2
X_10902_ _05750_ _02733_ _03371_ _03372_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11882_ _05033_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10833_ _00297_ _00810_ _00757_ _01365_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__nand4_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10764_ _03807_ _03808_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12503_ _05714_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10695_ _03731_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12434_ _05587_ _05640_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__xnor2_1
X_12365_ _05247_ _05258_ _05255_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__o21a_2
X_11316_ _04406_ _04414_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12296_ _05171_ _05151_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__and2b_1
X_11247_ _03817_ _03826_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__xnor2_1
X_11178_ _03768_ _03847_ _03845_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a21o_2
X_10129_ _02431_ _02436_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07340_ _00242_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09010_ _01908_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07271_ _00172_ _00173_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _02856_ _02873_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nand3_4
XFILLER_0_95_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09843_ net75 VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__buf_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _02046_ _02040_ _01412_ _02043_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__a2bb2o_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06297_ _06298_ _06252_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__a21oi_1
X_08725_ _01041_ _01602_ _01625_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__o21a_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _00059_ _00062_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__nand2_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _03260_ _00080_ _00507_ _02855_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22oi_1
X_08587_ net74 VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07538_ _02646_ _00438_ _00439_ _00440_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07469_ _05980_ _05969_ _00370_ _00371_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09208_ _02105_ _02106_ _01977_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__o21a_1
X_10480_ _05191_ net181 _03496_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09139_ _06375_ net10 VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12150_ _04956_ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11101_ _04178_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__or2b_2
XFILLER_0_130_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12081_ _05249_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11032_ _01002_ net196 VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__and2_1
X_11934_ _05076_ _05091_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11865_ _05003_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__xor2_1
X_10816_ _01293_ net146 _02615_ _06319_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11796_ _04547_ _04564_ _04941_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__a21o_1
X_10747_ _03778_ _03779_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10678_ _03713_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12417_ _05330_ _05332_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12348_ _01872_ _03210_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12279_ _05470_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__and2b_1
X_06840_ net121 _06151_ _06153_ _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__and4_1
X_06771_ _05805_ _05816_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__nor2_1
X_08510_ _03798_ _00850_ _01410_ _02470_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__a22o_1
X_09490_ _01731_ _01761_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21bo_1
X_08441_ _01339_ _01340_ _01286_ _00817_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08372_ _01262_ _01272_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07323_ _00225_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07254_ _06211_ _00156_ _00157_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07185_ _00087_ _00088_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09826_ _02764_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__xnor2_2
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ _02021_ _02023_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__nand2_1
X_06969_ net133 VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__clkbuf_4
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ net220 net229 net221 net228 VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__a22o_1
X_09688_ _06173_ net206 net207 _04106_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__a22o_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _01537_ _01538_ _01517_ _01518_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a211o_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _04306_ _04308_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10601_ _00109_ _00544_ net212 net223 VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__nand4_1
X_11581_ _04022_ _04219_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10532_ _02955_ _03554_ _02962_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10463_ _03464_ _03478_ _03476_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10394_ _03394_ _03402_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12202_ _05352_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12133_ _05306_ _04927_ _05309_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12064_ _04848_ _04877_ _05234_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11015_ _04082_ _04083_ _03506_ _03508_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11917_ _04647_ _04650_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__nand2_1
X_12897_ clknet_1_1__leaf_clk _00021_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dfxtp_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11848_ _04555_ _04997_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11779_ _04505_ _04506_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08990_ _01851_ _01852_ _01888_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__a211o_1
X_07941_ _00826_ _00841_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__nor2_1
X_07872_ net144 VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09611_ _01936_ _01952_ _01951_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__a21o_2
X_06823_ net17 VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09542_ net18 net29 net30 net17 VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a22o_1
X_06754_ _03469_ _05630_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nor2_1
X_06685_ _03084_ _02822_ _03194_ _04862_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__and4_1
X_09473_ _01727_ _02391_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__nand3_2
X_08424_ _04106_ _06172_ net204 net205 VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__nand4_1
X_08355_ net124 net125 _06283_ _00201_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__nand4_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07306_ net131 net125 net126 net130 VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08286_ _01186_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07237_ _00043_ _00139_ _00140_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__and3_2
X_07168_ _00057_ _00071_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07099_ _02668_ _06410_ _06411_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09809_ _02759_ _02760_ _02755_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a21o_1
X_12820_ _06006_ _06011_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ net264 _05900_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11702_ _04835_ _04837_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__xnor2_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05833_ _05835_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11633_ _04760_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11564_ _04198_ _04200_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10515_ _00480_ net187 net188 _00989_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__a22o_1
X_11495_ _04610_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nor2_1
X_10446_ _03453_ _03459_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10377_ _03335_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__xnor2_2
X_12116_ _04901_ _05291_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__nand2_1
X_12047_ _01264_ _01250_ _01872_ _03210_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06470_ _02470_ _02481_ _02492_ _02503_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__nand4_4
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08140_ _01035_ _01040_ _00511_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08071_ _00969_ _00972_ _00908_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07022_ _06301_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08973_ _04314_ _01264_ _01872_ net130 VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a22o_1
X_07924_ _00824_ _00825_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07855_ net214 VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__buf_2
X_07786_ _00663_ _00664_ _00687_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06806_ _06119_ _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__or2_1
X_06737_ net103 _05444_ _03535_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__nand3_1
X_09525_ _02412_ _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09456_ _02371_ _02373_ _01691_ _02198_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__a211o_1
X_06668_ _03042_ _04677_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__nand2_1
X_08407_ _00769_ _00770_ _00771_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06599_ net200 VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__clkbuf_4
X_09387_ _02296_ _02297_ _02267_ _01646_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08338_ _01237_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08269_ _00627_ _01168_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10300_ _03285_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11280_ _04374_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10231_ _03222_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10162_ _03146_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__xnor2_2
X_10093_ _03070_ _03071_ _03072_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12803_ net266 _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10995_ _03525_ _03529_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a21o_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _05966_ _05968_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _05891_ _05892_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__nand2_1
X_12596_ _01667_ _01652_ _03019_ _03006_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11616_ _04742_ _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__nor2_1
X_11547_ _04189_ _04197_ _04188_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11478_ _04565_ _04592_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__nor3_2
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10429_ _02817_ _03440_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ net37 VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07571_ _03381_ _00062_ _00472_ _00473_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__o2bb2a_1
X_06522_ net112 VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09310_ _02212_ _02213_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09241_ _01500_ _01502_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__nand2_1
X_06453_ _02317_ _02328_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09172_ net60 net61 net55 VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ net228 net220 net229 net219 VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ net108 VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_4
X_07005_ net151 VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput118 data_in[205] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xinput107 data_in[196] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput129 data_in[215] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_08956_ _04303_ net121 net137 net138 VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__and4_1
X_07907_ _00372_ _00373_ _00375_ _00376_ _00369_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a32o_1
X_08887_ net16 _06138_ _00647_ _01181_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__and4_1
X_07838_ _00314_ _00325_ _00739_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07769_ _00668_ _00669_ _00203_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09508_ _02428_ _02430_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10780_ _03823_ _03824_ _03825_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _02353_ _02354_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__and3_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _05650_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__xnor2_2
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11401_ net72 net84 VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12381_ _05518_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__xnor2_1
X_11332_ _04295_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11263_ net135 net136 net128 net129 VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10214_ _02567_ _02566_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__or2b_1
X_11194_ _04279_ _04280_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__nor2_1
X_10145_ _02479_ _02458_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10076_ _01764_ _02388_ _02387_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10978_ _03467_ _03470_ _03468_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__a21boi_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12717_ _05932_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12648_ _05874_ _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12579_ _05303_ _05592_ _05595_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _01708_ _01709_ _01173_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a21oi_2
X_09790_ _02035_ _02047_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__nor2_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _01634_ _01640_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__and3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _01570_ _01571_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07623_ _00506_ _00090_ _00525_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07554_ _00455_ _00456_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07485_ net52 _05761_ net53 _03743_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06505_ _02877_ _02888_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09224_ _02121_ _02122_ _01494_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09155_ _02003_ _02054_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09086_ net207 VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08106_ _00491_ _00493_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08037_ net69 net70 net80 net81 VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ net221 net230 VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__and2_1
X_08939_ _01836_ _01837_ net86 net101 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__and4bb_1
X_11950_ _04531_ _04704_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a21oi_2
X_10901_ _03943_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__xnor2_2
X_11881_ _01567_ _02239_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10832_ _00810_ net214 net206 _00297_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10763_ _03805_ _03806_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _05272_ _05465_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__a21boi_1
X_10694_ _03705_ _03706_ _03730_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12433_ _05589_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12364_ _05294_ _05317_ _05315_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11315_ _04406_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _05150_ _05172_ _05176_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__a21o_1
X_11246_ _03799_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nor2_1
X_11177_ _03731_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__nor2_2
X_10128_ _03109_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__or2_1
X_10059_ _02979_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__xor2_4
XFILLER_0_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07270_ _04227_ _06227_ _00171_ net157 VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09911_ _02871_ _02872_ _02857_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09842_ _06424_ _06410_ _00431_ _00421_ _02118_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__a41o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09773_ _02720_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__nor2_2
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _01065_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__xor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _06252_ _06297_ _06298_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08655_ _01554_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__nor2_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _00081_ _00508_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__nor2_1
X_08586_ net73 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07537_ _03524_ _05389_ _05444_ _06416_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__nand4_2
XFILLER_0_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07468_ net243 net244 net238 net239 VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__nand4_4
XFILLER_0_107_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07399_ net200 net211 _00299_ _00300_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__a22o_1
X_09207_ _01977_ _02105_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__nor3_1
XFILLER_0_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09138_ _02036_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11100_ _04168_ _03628_ _04177_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__or3_1
X_09069_ _01768_ _01769_ _01967_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12080_ _05251_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__and2_1
X_11031_ _00480_ net188 net189 _00989_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__a22o_1
X_11933_ _05076_ _05091_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11864_ _05006_ _05015_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__xnor2_1
X_10815_ _03863_ _03865_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11795_ _04561_ _04563_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10746_ _03788_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10677_ _03711_ _03712_ _01777_ _00617_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__and4bb_1
X_12416_ _04509_ _04510_ _04954_ _05327_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12347_ _05544_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12278_ _05467_ _05469_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__nand2_1
X_11229_ _00703_ net92 _01858_ _00238_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06770_ _02569_ _05750_ _05772_ _05794_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__a22oi_1
X_08440_ _01286_ _00817_ _01339_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_86_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ _01263_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07322_ _06136_ _06259_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07253_ _00154_ _00155_ _06225_ _06214_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07184_ _03227_ _02866_ _04741_ _00086_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09825_ _02777_ _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__xnor2_2
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _02693_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__xor2_2
X_06968_ _06273_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__xor2_4
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _02625_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__xor2_2
X_08707_ _03227_ _00516_ _01025_ _01026_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__and4_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _01517_ _01518_ _01537_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__o211ai_4
X_06899_ _06205_ _06206_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__or3_2
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08569_ net71 _06410_ _00421_ _05498_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__a22oi_1
X_10600_ net34 net212 net223 _00109_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a22o_1
X_11580_ _04215_ _04218_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10531_ _02960_ _02961_ _02956_ _02277_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10462_ _03461_ _03462_ _03463_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12201_ _05368_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10393_ _03400_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _05306_ _04927_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12063_ _04850_ _04876_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11014_ _03506_ _03508_ _04082_ _04083_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11916_ _05072_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12896_ clknet_1_1__leaf_clk _00020_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dfxtp_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11847_ _04557_ _04559_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__or2_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _04920_ _04921_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10729_ _00250_ _01217_ _02498_ _06264_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07940_ _00826_ _00841_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__and2_1
X_07871_ _00769_ _00770_ _00771_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__a21oi_1
X_09610_ _01871_ _01880_ _01881_ _01884_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__a31o_2
X_06822_ _06135_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09541_ _02465_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__or2_2
X_06753_ _05597_ _05608_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__and2_1
X_06684_ _03084_ _03194_ _04862_ _02822_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09472_ _02389_ _02390_ _01728_ _01710_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__a211o_1
X_08423_ _06172_ net204 net205 net209 VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08354_ net125 _06283_ _00201_ net124 VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07305_ _06279_ _06280_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08285_ net166 net162 net163 net165 VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07236_ _00137_ _00138_ _00044_ _05323_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o211ai_2
X_07167_ _00069_ _00070_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07098_ _02668_ _06410_ _06411_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__and3_1
X_09808_ _02755_ _02759_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__and3_1
X_09739_ _02683_ _02682_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__inv_2
X_11701_ _04346_ _04373_ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_84_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _05833_ _05835_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__nand2_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11632_ _04731_ _04732_ _04759_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11563_ _04685_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__nand2_2
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10514_ _00047_ net196 _02911_ _02912_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__and4_1
X_11494_ _00489_ _01002_ _01562_ _02904_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__and4_2
XFILLER_0_33_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10445_ _03456_ _03457_ _02859_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10376_ _03380_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__xnor2_2
X_12115_ _04901_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12046_ _01250_ _01872_ _03210_ _01264_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12879_ clknet_1_0__leaf_clk _00003_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dfxtp_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08070_ _00970_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07021_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08972_ net129 VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_4
X_07923_ _02481_ _00821_ _00823_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__a21oi_1
X_07854_ _00310_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06805_ _03996_ _06118_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07785_ _00323_ _00686_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06736_ net115 VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__clkbuf_4
X_09524_ _02414_ _02447_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__xnor2_4
X_09455_ _01691_ _02198_ _02371_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__o211ai_2
X_06667_ _03042_ _04677_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or2_1
X_08406_ _01305_ _01306_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09386_ _02267_ _01646_ _02296_ _02297_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06598_ _02525_ _03919_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__xnor2_1
X_08337_ _01228_ _00674_ _01236_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08268_ _00627_ _01168_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07219_ _02811_ _00107_ _00121_ _00122_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__nand4_2
XFILLER_0_116_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _03220_ _03221_ _03214_ _03215_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a211o_1
X_08199_ _00571_ net299 _01099_ _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__o211a_2
XFILLER_0_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10161_ _02471_ _02473_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__or2_1
X_10092_ _03070_ _03071_ _00166_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a21oi_1
X_10994_ _02906_ _03528_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__and2_1
X_12802_ _06040_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05766_ _05890_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__a21oi_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05891_ _05892_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11615_ _01188_ _01157_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__and2_1
X_12595_ _05679_ _05704_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11546_ _04661_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11477_ _04590_ _04591_ _04566_ _04082_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10428_ _00431_ net82 _03438_ _03439_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10359_ _02754_ _02762_ _02761_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _05195_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07570_ _03392_ _05191_ _05202_ _00059_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__and4_1
X_06521_ net33 VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09240_ _02131_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06452_ net157 VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09171_ _02068_ _02069_ _01446_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08122_ _02866_ _01023_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08053_ _03381_ net78 _00453_ _00953_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__nand4_2
X_07004_ _06182_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput108 data_in[197] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
X_08955_ _04303_ net137 net138 net121 VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__a22oi_1
Xinput119 data_in[206] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
X_07906_ _06371_ _00377_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08886_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__inv_2
X_07837_ _00290_ _00313_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__and2b_1
X_07768_ _00203_ _00668_ _00669_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06719_ _02734_ _05191_ _05213_ _05235_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__a22o_1
X_09507_ _01742_ _01743_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07699_ _00156_ _00168_ _00597_ _00598_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__o211ai_1
X_09438_ _01664_ _01674_ _01673_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _01610_ _01611_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__nand2_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ _03998_ _04003_ _04002_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_34_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12380_ _05521_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11331_ _04379_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_50_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11262_ net136 net128 net129 _00201_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_105_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10213_ _02566_ _02567_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__and2b_1
X_11193_ _04278_ _04268_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__and2b_1
X_10144_ _02667_ _02792_ _03127_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__a21o_2
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10075_ _02451_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10977_ _04042_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__or2_2
XFILLER_0_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12716_ _05933_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__xor2_2
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12647_ _05872_ _05873_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12578_ _05613_ _05614_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11529_ _04648_ _04649_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _01637_ _01638_ _01639_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__a21o_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08671_ _00988_ _00990_ _00991_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__a21bo_1
X_07622_ _00515_ _00524_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07553_ _02635_ _03546_ _06437_ _00454_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07484_ net54 VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06504_ _02778_ _02877_ _02888_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__and3_2
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09223_ _01494_ _02121_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09154_ _02052_ _02053_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08105_ _01005_ _01006_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__or2_1
X_09085_ _01384_ _01393_ _01392_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput90 data_in[180] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ net70 net80 net81 net69 VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09987_ net228 net229 net222 net224 VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nand4_1
X_08938_ net86 _01835_ _01836_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__o2bb2a_1
X_08869_ _01465_ _01357_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__or2b_1
X_10900_ _03957_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11880_ _00481_ _01584_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nand2_1
X_10831_ _03881_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10762_ _03805_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12501_ _05462_ _05464_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10693_ _03705_ _03706_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__a21oi_1
X_12432_ _05618_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12363_ _05240_ _05262_ _05260_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11314_ _04411_ _04412_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__xnor2_1
X_12294_ _05475_ _05148_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__or2b_1
X_11245_ _06134_ _01251_ _03212_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11176_ _03704_ _03734_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__and2b_1
X_10127_ _03107_ _03108_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__and2_1
X_10058_ _03033_ _03035_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09910_ _02857_ _02871_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__nand3_4
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09841_ _02131_ _02138_ _02137_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__a21bo_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _02718_ _02719_ _02704_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a21oi_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _06294_ _06296_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__nand2_1
X_08723_ _01616_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__xnor2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08654_ net174 net175 _00479_ _00985_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__and4_1
X_07605_ _02855_ _03260_ _00080_ _00507_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__nand4_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _03524_ net103 _00910_ _01484_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07536_ _05389_ _05444_ _06416_ _03524_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07467_ net244 net238 net239 net243 VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09206_ _02103_ _02104_ _01978_ _01979_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07398_ _03941_ _06304_ _00299_ _00300_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__nand4_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09137_ _05882_ _06368_ _00357_ _00850_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__nand4_1
XFILLER_0_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09068_ _01896_ _01897_ _01965_ _01966_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__a22oi_2
X_08019_ _05444_ _06437_ _06416_ _05389_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11030_ _00058_ _00481_ net188 net189 VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nand4_1
X_11932_ _05078_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11863_ _05013_ _05014_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__xnor2_1
X_10814_ _06311_ net155 VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11794_ _04497_ _04519_ _04938_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_131_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10745_ _06284_ net102 VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10676_ _01777_ _00617_ _03711_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12415_ _05325_ _05337_ _05335_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__a21oi_2
X_12346_ _05207_ _05217_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12277_ _05467_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__nor2_1
X_11228_ _04298_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__xnor2_1
X_11159_ net259 _04242_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08370_ _01269_ _01270_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ _00196_ _00223_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07252_ _06225_ _06214_ _00154_ _00155_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07183_ _03227_ _04741_ _00086_ _02866_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09824_ _02071_ _02076_ _02070_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__a21boi_2
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _02700_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__and2b_1
X_06967_ _06279_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__xor2_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ _06086_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__nand2_1
X_08706_ _04752_ _04741_ _00080_ _00086_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__and4_1
X_06898_ _06211_ _06212_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__nand2_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08637_ _01535_ _01536_ _01519_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__a21o_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _00939_ _00942_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08499_ _01398_ _01399_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__nand2_1
X_07519_ _03579_ _06410_ _00421_ _02668_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10530_ _02930_ _02936_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10461_ _03464_ _03465_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__and3b_1
X_12200_ _05382_ _05384_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10392_ _03398_ _03399_ _03395_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__a21o_1
X_12131_ _05307_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__xnor2_1
X_12062_ _05199_ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11013_ _04080_ _04081_ _03501_ _04059_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11915_ _04669_ _04670_ _04686_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__o21a_2
XFILLER_0_59_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12895_ clknet_1_1__leaf_clk _00019_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11846_ _04557_ _04559_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__and2_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04909_ _04919_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10728_ _00250_ _00706_ _03164_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__nand3_1
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10659_ _03124_ _03081_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12329_ _04775_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07870_ _00769_ _00770_ _00771_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__and3_1
X_06821_ _04292_ _02251_ _04424_ _06134_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__and4_1
X_09540_ _04238_ _06130_ _01188_ net164 VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__and4_1
X_06752_ _03469_ _05597_ _05608_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09471_ _01728_ _01710_ _02389_ _02390_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__o211ai_4
X_06683_ net43 VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__clkbuf_4
X_08422_ _06086_ _06304_ _00763_ _00764_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08353_ _01252_ _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07304_ _00205_ _00206_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__nand2_1
X_08284_ _01182_ _01184_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07235_ _00044_ _05323_ _00137_ _00138_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07166_ _00060_ _00061_ _00067_ _00068_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07097_ _05487_ _05531_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09807_ _05750_ _01434_ _02757_ _02758_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__nand4_2
X_07999_ net298 _00867_ _00899_ _00900_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__or4bb_1
X_09738_ _02682_ _02683_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09669_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__inv_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04370_ _04372_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__and2b_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05907_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__xor2_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _04731_ _04732_ _04759_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a21oi_1
X_11562_ _04671_ _04684_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10513_ _00058_ _00489_ _00481_ _01002_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11493_ _01002_ _01562_ _02904_ _00489_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10444_ _02859_ _03456_ _03457_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10375_ _02722_ _02743_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12114_ _05288_ _05289_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12045_ _04854_ _04857_ _04858_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12878_ clknet_1_0__leaf_clk _00002_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dfxtp_2
X_11829_ _04540_ _04541_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07020_ _06189_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08971_ _01270_ _01269_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07922_ _02481_ _00821_ _00823_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__and3_1
X_07853_ _00320_ _00754_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__xnor2_2
X_06804_ _03996_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__nor2_1
X_07784_ _00676_ _00685_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__xnor2_1
X_06735_ _03425_ _05422_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__xnor2_1
X_09523_ _02416_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__xnor2_4
X_09454_ _02369_ _02370_ _02264_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__a21o_1
X_06666_ net269 _04666_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__xnor2_1
X_08405_ _01303_ _01304_ _01287_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__a21o_1
X_09385_ _02293_ _02294_ _02281_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06597_ _03842_ _03908_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__xor2_4
X_08336_ _01228_ _00674_ _01236_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08267_ _01140_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07218_ _00119_ _00120_ _00108_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08198_ _01097_ _01098_ _01046_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07149_ _05126_ _05147_ _00051_ _00052_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__a211o_1
X_10160_ _03144_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__xnor2_2
X_10091_ _02403_ _02406_ _02402_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10993_ _03496_ _03500_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__nand2_1
X_12801_ _06041_ _05982_ _05975_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__o21a_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _05887_ _05889_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__nor2_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05516_ _05719_ _05717_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11614_ _04273_ _04740_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__xor2_1
X_12594_ _05676_ _05678_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11545_ _04193_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11476_ _04566_ _04082_ _04590_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__a211oi_2
X_10427_ _00431_ net82 _03438_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10358_ _02728_ _02729_ _02737_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _03286_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12028_ _04783_ _05185_ _05194_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06520_ _02437_ _02987_ _02998_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06451_ net165 VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09170_ _01446_ _02068_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08121_ net231 VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08052_ net89 _00453_ _00953_ net78 VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07003_ _06310_ _06316_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput109 data_in[198] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_4
X_08954_ _01262_ _01272_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07905_ _00345_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__inv_2
X_08885_ net17 net29 net30 net16 VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__a22o_1
X_07836_ _00383_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07767_ net121 _00665_ _00666_ _00667_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__nand4_2
X_06718_ _02734_ _05191_ _05213_ _05235_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nand4_2
X_09506_ _01736_ _01741_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07698_ _00160_ _00599_ _00600_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__or3b_1
X_09437_ _02351_ _02352_ _02343_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06649_ _02251_ _04424_ _04457_ _04479_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ _02276_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08319_ _02196_ _04446_ _00706_ _01217_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__and4_1
X_09299_ _00059_ _00062_ _01556_ _01555_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11330_ _04429_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11261_ _04352_ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__and2_1
X_10212_ _03187_ _03202_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__xnor2_1
X_11192_ _04268_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__and2b_1
X_10143_ _02791_ _02669_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10074_ _03051_ _03052_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ _04038_ _04039_ _04041_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12715_ _05935_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12646_ _05872_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12577_ _05566_ _05573_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11528_ _00543_ _04154_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11459_ _00985_ _01524_ _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ net183 _01567_ _01568_ _01569_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__a22o_1
X_07621_ _00522_ _00523_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__nand2_1
X_07552_ _03546_ _06437_ _00454_ _02635_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06503_ _02833_ _02844_ _02855_ _02866_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07483_ _06348_ _06350_ _02569_ _06343_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__and4b_1
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09222_ _02119_ _02120_ _02114_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09153_ _01403_ _01423_ _01421_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08104_ _01003_ _01004_ net193 _00049_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09084_ _01395_ _01982_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput91 data_in[181] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput80 data_in[171] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08035_ net82 VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09986_ net229 net222 net224 net228 VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__a22o_1
X_08937_ net87 net88 net98 net99 VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__and4_1
X_08868_ _01358_ _01464_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07819_ _00719_ _00720_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__nor2_1
X_08799_ _01105_ _01107_ _01697_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o211ai_4
X_10830_ _03287_ _03879_ _03880_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10761_ _03188_ _03198_ _03197_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10692_ _03728_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__xor2_1
X_12500_ _05583_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12431_ _05636_ _05637_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12362_ _05539_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11313_ _03887_ _03888_ _03891_ _03292_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12293_ _05473_ _05474_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__or2_1
X_11244_ _03797_ _03801_ _03803_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ _03740_ _03914_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a21o_2
X_10126_ _03107_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__nor2_1
X_10057_ _02325_ _02362_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10959_ _03523_ _03566_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12629_ _05681_ _05703_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09840_ _02119_ _02121_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand2_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09771_ _02704_ _02718_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__and3_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _06294_ _06296_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08722_ _01037_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__xnor2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _05202_ _00479_ _00985_ _03392_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07604_ net221 VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__buf_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08584_ _03524_ _00910_ _01484_ _02646_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_119_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07535_ net117 VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_4
X_07466_ _00367_ _00368_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ _01978_ _01979_ _02103_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07397_ _06077_ net210 net203 net209 VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09136_ _06368_ net2 _00850_ _05882_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09067_ _01896_ _01897_ _01965_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__and4_1
X_08018_ _00440_ _00441_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__nand2_1
X_09969_ _02929_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__xor2_2
X_11931_ _05084_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11862_ _04577_ _04580_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10813_ net153 _03861_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11793_ _04499_ _04518_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10744_ _03785_ _03786_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10675_ _06227_ net164 _03709_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12414_ _05320_ _05341_ _05339_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12345_ _04795_ _05541_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12276_ _04889_ _05112_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11227_ _04299_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__xor2_1
X_11158_ net259 _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__nand2_1
X_10109_ _02438_ _02439_ _02443_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__o21ba_2
X_11089_ _03611_ _03613_ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__a21o_2
XFILLER_0_78_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07320_ _00221_ _00222_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07251_ _00152_ _00153_ _06241_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a21oi_2
X_07182_ net229 VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09823_ _02771_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _02698_ _02699_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__or2_1
X_06966_ net121 _06151_ _06154_ _04336_ _06152_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a32o_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09685_ net215 VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__buf_2
X_08705_ _01604_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__nor2_1
X_06897_ _06210_ _06207_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__or2b_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _01519_ _01535_ _01536_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__nand3_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08567_ _00526_ _01017_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__and2_1
X_08498_ _03820_ net252 _00821_ _01397_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__nand4_1
XFILLER_0_91_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07518_ net81 VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__buf_2
X_07449_ _00350_ _00351_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10460_ _03466_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09119_ net14 VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10391_ _03395_ _03398_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12130_ _01444_ _03967_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12061_ _05229_ _05231_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11012_ _03501_ _04059_ _04080_ _04081_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a211o_2
XFILLER_0_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11914_ _05063_ _05070_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12894_ clknet_1_1__leaf_clk _00018_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfxtp_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11845_ _04993_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__nand2_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _04909_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10727_ _03237_ _03240_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10658_ _03123_ _03082_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10589_ _03616_ _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__or2b_2
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12328_ _02498_ _01784_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12259_ _05432_ _05092_ _05448_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__or3_1
X_06820_ _04292_ _04424_ _06134_ _02251_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__a22oi_1
X_06751_ _05433_ _05586_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06682_ _04818_ _04840_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__nor2_1
X_09470_ _02387_ _02388_ _01764_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__a21o_1
X_08421_ _04106_ _06173_ _06362_ _00343_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08352_ net121 net94 _01250_ _01251_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__and4_2
XFILLER_0_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07303_ _02240_ _00200_ _00202_ _00204_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08283_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07234_ _00135_ _00136_ _00077_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07165_ _00060_ _00061_ _00067_ _00068_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__nor4_1
XFILLER_0_14_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07096_ net80 VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09806_ _05750_ net65 _02757_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__a22o_1
X_07998_ _00897_ _00898_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09737_ _02030_ _02028_ _02032_ _02018_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__a22o_1
X_06949_ net24 net25 _06138_ _06261_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09668_ _02604_ _02605_ _02587_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09599_ _02529_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__nand2_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08619_ net109 VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_4
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11630_ _04734_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11561_ _04671_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10512_ _03531_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nor2_1
X_11492_ _04607_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10443_ _00438_ _00956_ _03454_ _03455_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nand4_1
X_10374_ _02742_ _02740_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__and2b_1
X_12113_ _05277_ _04921_ _05287_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12044_ _04365_ _04830_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12877_ clknet_1_0__leaf_clk _00001_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dfxtp_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _04603_ _04632_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11759_ _04445_ _04449_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08970_ _01868_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__nor2_1
X_07921_ _02481_ _00822_ _00351_ _00350_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__a31o_1
X_07852_ _00752_ _00753_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__and2b_1
Xinput1 data_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_06803_ _06116_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__or2_1
X_07783_ _00215_ _00684_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09522_ _02417_ _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__xor2_4
X_06734_ _05400_ _05411_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__or2_1
X_09453_ _02264_ _02369_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__nand3_1
X_06665_ _02350_ _04655_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__xor2_2
X_08404_ _01287_ _01303_ _01304_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__nand3_4
X_09384_ _02281_ _02293_ _02294_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__and3_1
X_06596_ _03875_ _03897_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nand2_2
X_08335_ _01234_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08266_ _01141_ _01166_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07217_ _00108_ net317 _00120_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08197_ _01046_ _01097_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07148_ _03337_ _05093_ _00048_ _00050_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07079_ _02503_ _06383_ _06391_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10090_ _03069_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12800_ _05977_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__inv_2
X_10992_ _03530_ _03549_ _03548_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _05954_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _05766_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _03709_ _02464_ _00617_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ _05768_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11544_ _04662_ _04665_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11475_ _04587_ _04588_ _04568_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10426_ _06410_ net81 net73 net74 VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10357_ _02732_ _02733_ _02736_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _00343_ net213 net205 net214 VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__and4_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ _04783_ _05185_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06450_ _02196_ _02207_ _02262_ _02284_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08120_ _01021_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08051_ net178 VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_4
X_07002_ _06313_ _06314_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _01263_ _01271_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__or2_1
X_07904_ _00805_ _00408_ _00412_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08884_ net31 VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07835_ _00734_ _00735_ _00659_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__o21a_1
X_07766_ net121 _00665_ _00666_ _00667_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06717_ _05224_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09505_ _02425_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__xor2_1
X_09436_ _02343_ _02351_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07697_ _00597_ _00598_ _00156_ _00168_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__a211o_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06648_ _02207_ _04468_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__nand2_1
X_09367_ _00080_ net230 _02274_ _02275_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__and4_2
X_06579_ _03689_ _03699_ _02943_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09298_ _01065_ _01624_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__nor2_1
X_08318_ _01218_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08249_ _01143_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11260_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10211_ _03200_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__xor2_1
X_11191_ _04276_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__xnor2_1
X_10142_ _02659_ _02661_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10073_ _01973_ _02384_ _02382_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10975_ _04038_ _04039_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__a21oi_1
X_12714_ _05938_ _05946_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__xor2_2
XFILLER_0_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12645_ _05621_ _05633_ _05632_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__o21ba_1
X_12576_ _05288_ _05293_ _05572_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11527_ _00543_ _01629_ _04171_ _04170_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11458_ _00453_ _00953_ _01563_ _02215_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nand4_2
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10409_ _03391_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__xnor2_2
X_11389_ _04004_ _04006_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07620_ _00088_ _00521_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07551_ net107 VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_4
X_06502_ _02833_ _02844_ _02855_ _02866_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07482_ _06415_ _06431_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09221_ _02114_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09152_ _02033_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08103_ _05093_ _00049_ _01003_ _01004_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__o2bb2a_1
X_09083_ _00824_ _01401_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput81 data_in[172] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput70 data_in[162] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
XFILLER_0_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08034_ _00932_ _00933_ _00934_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput92 data_in[182] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09985_ _04741_ _00086_ _00507_ _01034_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__and4_1
X_08936_ net88 _00238_ _00703_ net87 VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__a22oi_1
X_08867_ _01349_ _01351_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__and2b_1
X_07818_ _06159_ net97 _00717_ _00718_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _01549_ _01550_ _01698_ _01696_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07749_ _00252_ _00641_ _00650_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__o21ai_2
X_10760_ _03803_ _03804_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__nand2_1
X_09419_ _02327_ _02332_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10691_ _06243_ net173 VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12430_ _05635_ _05620_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12361_ _05559_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11312_ _04409_ _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__xnor2_1
X_12292_ _05483_ _05484_ _05485_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11243_ _04332_ _04334_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__xnor2_2
X_11174_ _03913_ _03741_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__and2b_1
X_10125_ _06243_ net172 VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__and2_1
X_10056_ _02326_ _01680_ _02358_ _02359_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10958_ _03510_ _03512_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__or2b_2
XFILLER_0_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10889_ net3 net11 net13 net2 VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12628_ _05682_ _05702_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12559_ _05773_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09770_ _02714_ _02715_ _02717_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _04391_ _06161_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__o21a_1
X_08721_ _01620_ _01621_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__and2b_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _05191_ _00062_ _00979_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__and3_1
X_07603_ _04796_ _00084_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08583_ net119 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07534_ _00436_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__inv_2
X_07465_ _03853_ net235 _06383_ _00366_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09204_ _02101_ _02102_ _02055_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07396_ net209 _06077_ _06172_ _06361_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__nand4_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09135_ _00874_ _01440_ _01439_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09066_ _01963_ _01964_ _01345_ _01898_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__a211o_1
X_08017_ _00917_ _00918_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09968_ _02930_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08919_ _01203_ _01205_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__nand2_1
X_11930_ _05085_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__xor2_1
X_09899_ net100 _00059_ _00453_ _00953_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__and4_1
X_11861_ _05011_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__xor2_2
X_10812_ net144 net153 net154 net143 VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__a22o_1
X_11792_ _04908_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10743_ _03174_ _03176_ _03784_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__nor3_1
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10674_ _06227_ _02464_ _03709_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ _05616_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__or2b_2
XFILLER_0_63_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12344_ _01251_ _01835_ _01858_ _03180_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__and4_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12275_ _05109_ _05111_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__nor2_1
X_11226_ _04301_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11157_ _04236_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10108_ _03087_ _02577_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__o21a_2
X_11088_ _03608_ _03614_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__and2b_1
X_10039_ net201 net34 net212 net23 VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07250_ _06241_ _00152_ _00153_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__and3_2
X_07181_ _04796_ _00084_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09822_ _02774_ _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__xor2_1
X_09753_ _02698_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__and2_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06277_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__xor2_4
X_08704_ _03227_ net217 _01023_ _01603_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__and4_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09684_ _00297_ _02622_ _02623_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__a21bo_1
X_06896_ _06207_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__or2b_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _00959_ _01533_ _01534_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__nand3_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ net307 _00460_ _00965_ _00967_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07517_ _06423_ _06425_ _03579_ _05520_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08497_ _03820_ _00821_ _01397_ net252 VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07448_ net254 net8 net9 net253 VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ _00266_ _00280_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__and2_1
X_09118_ _02008_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__xor2_4
XFILLER_0_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10390_ _06343_ net65 _03396_ _03397_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__nand4_2
X_09049_ _01942_ _01947_ _01948_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12060_ _04814_ _04834_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__o21ba_2
X_11011_ _04078_ _04079_ _04060_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a21oi_1
X_11913_ _05066_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__xor2_4
X_12893_ clknet_1_1__leaf_clk _00017_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11844_ _04048_ _04992_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or2_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _04916_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _03744_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10657_ _03070_ _03071_ _03686_ _03067_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__a211o_1
X_10588_ _03603_ _03011_ _03615_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12327_ _05187_ _05188_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12258_ _05432_ _05092_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o21ai_2
X_11209_ _04296_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__nand2_1
X_12189_ _00953_ _01563_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06750_ _05433_ _05586_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__or2_1
X_06681_ _02866_ _04741_ _04829_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a21oi_1
X_08420_ _01319_ _01320_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08351_ _02229_ _01250_ _01251_ net94 VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07302_ _02240_ _00200_ _00202_ _00204_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__nand4_2
X_08282_ net16 net15 net29 _01181_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__and4_1
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07233_ _00077_ _00135_ _00136_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__nor3_2
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07164_ _00065_ _00066_ _05224_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07095_ _05290_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09805_ net53 net54 _00397_ _00872_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__nand4_2
X_07997_ _00897_ _00898_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__or2_1
X_09736_ _02671_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__xnor2_1
X_06948_ _04446_ _06138_ _06261_ _02196_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__a22oi_2
X_09667_ _02587_ _02604_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__and3_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _00984_ _00999_ _00998_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__o21bai_2
X_06879_ _06192_ _06193_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__and2_1
X_09598_ _02527_ _02528_ _02523_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__a21o_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _05761_ net54 net55 _03743_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__a22o_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11560_ _04673_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10511_ _05115_ _00049_ net197 net198 VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__and4_2
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11491_ _04103_ _04104_ _04102_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10442_ net117 net108 _03454_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10373_ _03362_ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12112_ _05277_ _04921_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12043_ _05206_ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12876_ clknet_1_0__leaf_clk _00000_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dfxtp_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _04604_ _04631_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__or2b_1
XFILLER_0_68_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _04443_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10709_ _03146_ _03147_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__and2b_1
X_11689_ _04816_ _04822_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ net10 VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07851_ _00750_ _00751_ _00295_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__a21o_1
Xinput2 data_in[100] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_07782_ _00682_ _00683_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__xnor2_1
X_06802_ _03656_ _06115_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06733_ net104 net113 net114 _05389_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__and4_1
X_09521_ _02418_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__xor2_4
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _02367_ _02368_ _01686_ net311 VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__o211ai_4
X_06664_ _03073_ _04644_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__xnor2_2
X_08403_ _01301_ _01302_ _00778_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__a21o_1
X_09383_ _02290_ _02291_ _02292_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__a21o_1
X_06595_ _02503_ _03886_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08334_ _01232_ _01233_ _01229_ _00720_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_59_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08265_ _01164_ _01165_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07216_ net315 _00118_ _00110_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08196_ net301 _01096_ _01047_ _01048_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07147_ _03337_ _05093_ _00048_ _00050_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_15_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07078_ _02503_ _06383_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09719_ _02105_ _02107_ _02661_ _02662_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__o211a_1
X_10991_ _03487_ _03501_ _03503_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _05955_ _05964_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _05887_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _04298_ _04318_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__and2_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12592_ _05770_ _05813_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__xnor2_1
X_11543_ _04663_ _04664_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11474_ _04568_ _04587_ _04588_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__nor3_1
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10425_ net81 net73 net74 net80 VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10356_ _03345_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__xnor2_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _00297_ _00810_ _00757_ _00343_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _05192_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12859_ _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08050_ _00478_ _00487_ _00951_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__o21ai_1
X_07001_ _06178_ _04150_ _06312_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08952_ _01274_ _01248_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__or2b_1
X_07903_ _06359_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__inv_2
X_08883_ _01781_ _01782_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__nor2_1
X_07834_ _00659_ _00734_ _00735_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__nor3_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07765_ net122 net124 net133 net135 VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__nand4_2
XFILLER_0_79_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06716_ net89 _03392_ net78 _05202_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and4_1
X_07696_ _00156_ _00168_ _00597_ _00598_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__o211a_1
X_09504_ _01737_ _01740_ _01738_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o21ba_1
X_09435_ _02347_ _02348_ _02349_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06647_ _04435_ _02196_ _04446_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _00080_ _00516_ _02274_ _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06578_ _02943_ _03689_ _03699_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09297_ _01581_ _01595_ _02199_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__o21a_1
X_08317_ _04446_ _00706_ _01217_ _02196_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08248_ _01147_ _01148_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08179_ _01078_ _01079_ _01080_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10210_ _02520_ _02534_ _02533_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__o21ba_1
X_11190_ _01777_ _01157_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10141_ _03081_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__xnor2_2
X_10072_ _02666_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10974_ _06437_ _02132_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__and2_1
X_12713_ _05944_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12644_ _05869_ _05870_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12575_ _05793_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11526_ _00107_ _04154_ _04153_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11457_ _00953_ net145 _02215_ _00453_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__a22o_1
X_10408_ _03393_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__xnor2_2
X_11388_ _04037_ _04057_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__a21o_1
X_10339_ _03864_ _02694_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _04736_ _04756_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a21o_2
XFILLER_0_108_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07550_ net177 VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06501_ net217 VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__buf_2
XFILLER_0_124_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07481_ _00381_ _00382_ _00348_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09220_ _02117_ _02118_ _01490_ _01492_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_29_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09151_ _02049_ _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09082_ _01402_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08102_ net191 net192 net186 net187 VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08033_ _00932_ _00933_ _00934_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput71 data_in[163] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xinput82 data_in[173] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
Xinput60 data_in[153] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_0_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput93 data_in[183] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09984_ _02952_ _02953_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__xnor2_2
X_08935_ net101 VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08866_ _01355_ _01356_ _01704_ _01705_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__and4_1
X_07817_ _06159_ _06253_ _00717_ _00718_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a22oi_1
X_08797_ _01101_ net323 _01693_ _01694_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__o211ai_1
X_07748_ _00648_ _00649_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07679_ _00470_ _00471_ _00579_ _00580_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__a2bb2o_2
X_09418_ net41 _02329_ _02330_ _02331_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__nand4_1
XFILLER_0_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10690_ _03726_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09349_ _02233_ _02234_ _02255_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_105_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12360_ _05226_ _05540_ _05558_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nor3_1
XFILLER_0_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11311_ _00810_ _02626_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12291_ _05483_ _05484_ _02185_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11242_ _00250_ _02498_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ _03702_ _03736_ _04257_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__a21bo_2
X_10124_ _03104_ _03105_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ _03002_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10957_ _03917_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__xor2_4
XFILLER_0_128_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10888_ _03366_ _03369_ _03367_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_128_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12627_ _05618_ _05637_ _05636_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_81_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12558_ _05775_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__and2_1
X_11509_ _04625_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12489_ _05688_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _06150_ _06163_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08720_ _01618_ _01619_ _01053_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__a21o_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _01022_ _01045_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__o21a_1
X_07602_ _00131_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__inv_2
X_08582_ _01478_ _01479_ _01481_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__o21ai_2
X_07533_ _00434_ _00435_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07464_ _03853_ _06383_ _00366_ _02503_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09203_ _02055_ _02101_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09134_ _01404_ _01412_ _01414_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__o21bai_4
X_07395_ _02459_ _00297_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09065_ _01345_ _01898_ _01963_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__o211ai_4
X_08016_ _00911_ _00916_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09967_ _02931_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__xor2_2
X_08918_ _01237_ _01804_ _01816_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__nor3_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _02858_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__nor2_2
X_08849_ _01747_ _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__nor2_1
X_11860_ _00985_ _03499_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__nand2_1
X_10811_ net143 net144 net154 VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__and3_1
X_11791_ _04933_ _04935_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10742_ _03174_ _03176_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10673_ net170 _01188_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__and2_1
X_12412_ _05596_ _05615_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _01858_ _03180_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ _05272_ _05465_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11225_ _04302_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11156_ _03065_ _04237_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__a21o_1
X_11087_ _04138_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__xor2_4
X_10107_ _02575_ _02576_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__or2b_1
Xinput250 data_in[94] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_2
X_10038_ net23 net201 net34 VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11989_ _04746_ _04748_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07180_ _04785_ _00081_ _00083_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09821_ _02065_ _02067_ _02066_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__a21bo_1
X_09752_ _02009_ _02011_ _02010_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__a21bo_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _04303_ net132 VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__and2_2
X_08703_ _03227_ _01023_ _01603_ net217 VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__a22oi_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09683_ net204 net213 net214 _06361_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__a22o_1
X_06895_ _04281_ _04578_ _06208_ _06209_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _01533_ _01534_ _00959_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__a21o_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08565_ _01357_ _01465_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07516_ _00139_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08496_ net13 VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07447_ net253 net254 net8 net9 VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07378_ _00266_ _00280_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09117_ _02015_ _02016_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _01945_ _01946_ _01296_ _01298_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_115_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11010_ _04060_ _04078_ _04079_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11912_ _05067_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__nor2_2
X_12892_ clknet_1_1__leaf_clk _00016_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfxtp_1
X_11843_ _04048_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__nand2_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04465_ _04466_ _04464_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10725_ _03746_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10656_ _03685_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10587_ _03603_ _03011_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12326_ _05205_ _05200_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12257_ _05443_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11208_ _03747_ _03764_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__or2b_1
X_12188_ _00985_ _03499_ _05011_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__a31o_1
X_11139_ _03431_ _03665_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__a21oi_4
X_06680_ _04774_ _04785_ _04807_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08350_ net92 VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07301_ _00203_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08281_ _04435_ _00647_ _01181_ net15 VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07232_ _00133_ _00134_ _00078_ _00079_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07163_ _05224_ _00065_ _00066_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _05356_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09804_ net54 net63 net64 net53 VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07996_ _06357_ _00407_ _00406_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__a21o_1
X_09735_ _02672_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06947_ net18 VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__clkbuf_4
X_09666_ _02601_ _02603_ _02594_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__a21o_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _00458_ _00962_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__and2_1
X_06878_ _06169_ _06191_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__or2_1
X_09597_ _02523_ _02527_ _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__nand3_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _03743_ _05761_ net54 VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__and3_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08479_ _06384_ _06383_ _00366_ _05980_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11490_ _04605_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__nor2_1
X_10510_ _00049_ _01562_ _02904_ _05115_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10441_ net115 net116 net109 net110 VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nand4_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10372_ _03376_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__xor2_2
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12111_ _05285_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12042_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12875_ _06111_ _06113_ _00166_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a21oi_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11826_ _04592_ _04594_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _04458_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10708_ _03170_ _03186_ _03184_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11688_ _04819_ _04820_ _04821_ _04817_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10639_ _02666_ _03050_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12309_ _05499_ _05500_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__a21oi_1
X_07850_ _00295_ _00750_ _00751_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__and3_1
X_07781_ _02218_ _04314_ _06274_ _00210_ _00213_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a41o_1
X_06801_ _03656_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__and2_1
Xinput3 data_in[101] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
X_06732_ _03524_ _03546_ _05389_ _02635_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__a22oi_1
X_09520_ _02442_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09451_ _01686_ _01688_ _02367_ _02368_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__a211o_1
X_06663_ _04622_ _04633_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__nand2_1
X_08402_ _00778_ _01301_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__nand3_4
X_06594_ net236 net243 net244 VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__and3_1
X_09382_ _02290_ _02291_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nand3_1
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ _01229_ _00720_ _01232_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08264_ _01142_ _00657_ _01163_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07215_ _00110_ _00117_ _00118_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__or3_4
X_08195_ _01047_ _01048_ net301 _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_104_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07146_ _02712_ _03348_ _05115_ _00049_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__nand4_1
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07077_ _06389_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07979_ _05761_ net53 _00387_ _03743_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__a22o_1
X_09718_ _02659_ _02660_ _02578_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__a21o_1
X_10990_ _04037_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__xnor2_4
X_09649_ _01947_ _01949_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05583_ _05713_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11611_ _04299_ _04317_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__and2_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12591_ _05796_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__xnor2_1
X_11542_ _00550_ _01666_ net56 _03006_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__and4_2
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11473_ _04585_ _04586_ _04569_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10424_ _02803_ _02805_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10355_ _03358_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__or2b_2
XFILLER_0_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _03283_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ _04803_ _05190_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12858_ _06092_ _06097_ _06090_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__or3_4
XFILLER_0_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11809_ _04511_ _04954_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12789_ _06026_ _06028_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07000_ _04139_ _06178_ _06311_ _02383_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08951_ _01249_ _01273_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08882_ _01780_ _01777_ net168 _01778_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__and4b_1
X_07902_ _00418_ _00583_ net312 VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__or3_2
X_07833_ _00660_ _00661_ _00733_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__and3_1
X_07764_ net124 net133 net135 net122 VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06715_ _03381_ _03392_ _02745_ _05202_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07695_ _00595_ _00596_ _06236_ _06240_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__a211o_1
X_09503_ _02419_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__xnor2_1
X_09434_ _02347_ _02348_ _02349_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__nand3_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06646_ _04435_ _02196_ _04446_ _02207_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09365_ net228 net229 net221 net222 VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__nand4_1
X_06577_ _03513_ _03678_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08316_ net21 VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__buf_2
X_09296_ _01593_ _01594_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08247_ net158 _00617_ _01146_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08178_ net256 net201 net212 _02789_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07129_ _00031_ _00032_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10140_ _03082_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__xor2_2
X_10071_ _03048_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__xor2_4
X_10973_ _00454_ _00956_ _00910_ _01484_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__nand4_1
X_12712_ _05803_ _05939_ _05943_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12643_ _05866_ _05868_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ _05781_ _05792_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11525_ _04642_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11456_ _04071_ _04075_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10407_ _03404_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__xor2_2
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11387_ _04056_ _04055_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10338_ _03340_ _03341_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nand2_2
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _03263_ _03264_ _03265_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12008_ _04757_ _04735_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07480_ _00348_ _00381_ _00382_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__and3_2
X_06500_ net226 VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09150_ _01416_ _01418_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09081_ _00811_ _01373_ _01980_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__o21a_1
X_08101_ net192 _00489_ _01002_ net191 VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_114_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08032_ _06419_ _00443_ _00444_ _00448_ _00437_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput72 data_in[164] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
Xinput50 data_in[144] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput61 data_in[154] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
Xinput94 data_in[184] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
Xinput83 data_in[174] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09983_ net218 net233 VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08934_ _01833_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08865_ _01704_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__inv_2
X_07816_ _04413_ _06254_ net88 net90 VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__nand4_1
X_08796_ _01549_ _01550_ _01695_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__or4b_4
XFILLER_0_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07747_ _00645_ _00646_ _02207_ _00647_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07678_ _00470_ _00471_ _00579_ _00580_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__or4bb_4
X_09417_ net41 _02329_ _02330_ _02331_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06629_ _02328_ _04259_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09348_ _02250_ _02252_ _02254_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__a21o_1
X_11310_ _04407_ _04408_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09279_ _02177_ _02178_ _01559_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12290_ _05138_ _05142_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11241_ _06264_ _01217_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11172_ _03703_ _03735_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10123_ _03093_ _03094_ _03103_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10054_ _03029_ _03030_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10956_ _04019_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10887_ _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12626_ _05850_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12557_ _05543_ _05774_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11508_ _04126_ _04129_ _04626_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12488_ _05699_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11439_ _00454_ _02132_ _04548_ _04549_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__nand4_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06980_ _06292_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _00540_ _01044_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07601_ _00502_ _00503_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08581_ _01478_ _01479_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__or3_4
XFILLER_0_44_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07532_ _05498_ net79 _00432_ _00433_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__nand4_1
X_07463_ net248 VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09202_ _02099_ _02100_ _02056_ _02057_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07394_ net213 VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__buf_2
X_09133_ _02018_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__xor2_4
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09064_ _01961_ _01962_ _01899_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08015_ _00911_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09966_ _02933_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__xor2_2
X_08917_ _01237_ _01804_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__o21a_1
X_09897_ net89 net114 net181 net110 VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__and4_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _04227_ _01157_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__and2_1
X_08779_ _01659_ _01678_ _01679_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__and3_2
X_10810_ _06086_ _03859_ _03279_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11790_ _04474_ _04485_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o21a_1
X_10741_ _03782_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12411_ _05596_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__nor2_1
X_10672_ _03101_ _03102_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12342_ _05212_ _05228_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12273_ _05462_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11224_ _03759_ _04313_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__xnor2_1
X_11155_ _03074_ _04239_ _03682_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__a21oi_1
X_11086_ _04162_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__nor2_2
X_10106_ _02484_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__inv_2
Xinput251 data_in[95] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
Xinput240 data_in[85] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_2
X_10037_ _03011_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11988_ _04835_ _04837_ _04839_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_85_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10939_ _03409_ _03999_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12609_ _05831_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09820_ _02772_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nor2_1
X_09751_ _02696_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__nor2_1
X_06963_ _06275_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nand2_2
X_08702_ net232 VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__buf_2
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _06361_ _00343_ net214 VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__and3_1
X_06894_ _04270_ _04556_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__or2_1
X_08633_ _01531_ _01532_ _00982_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__a21o_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08564_ _01358_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07515_ _00416_ _00417_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__or2_1
X_08495_ _00845_ _00847_ _00846_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__a21bo_1
X_07446_ _06382_ _06394_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07377_ _00268_ _00279_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09116_ _02012_ _02013_ _02014_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09047_ _01296_ _01298_ _01945_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09949_ _02913_ _02914_ _02908_ _02909_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a211o_1
X_11911_ _01051_ _01653_ _01629_ _02329_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__and4_1
X_12891_ clknet_1_0__leaf_clk _00015_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dfxtp_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11842_ _04990_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__xnor2_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _04914_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__xor2_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _03747_ _03764_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10655_ _03687_ _03688_ _03690_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10586_ _03608_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__xnor2_1
X_12325_ _05206_ _05211_ _04808_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _05445_ _05446_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11207_ _03748_ _03763_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__or2b_1
X_12187_ _05007_ _05008_ _05010_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__and3_1
X_11138_ _03662_ _03664_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nor2_1
X_11069_ _04143_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07300_ net122 net121 _06283_ _00201_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08280_ net30 VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__buf_2
XFILLER_0_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07231_ _00078_ _00079_ _00133_ _00134_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__o211a_2
XFILLER_0_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07162_ _02745_ _00062_ _00063_ _00064_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07093_ _06404_ _06405_ _06112_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09803_ _06347_ _00387_ _02073_ _02072_ _01444_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__a32o_1
X_07995_ _00403_ _00896_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__xnor2_1
X_09734_ _02673_ _02678_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__xnor2_1
X_06946_ _06136_ _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__xnor2_1
X_09665_ _02594_ _02601_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__nand3_1
X_06877_ _06169_ _06191_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__nand2_1
X_08616_ _00959_ _00960_ _00476_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__and3b_1
X_09596_ net97 _00672_ _02524_ _02526_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__nand4_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _06343_ _06347_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__nand2_1
X_08478_ _00844_ _00860_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07429_ _06329_ _06328_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__and2b_2
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10440_ net116 net109 net110 net115 VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10371_ _02724_ _02739_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12110_ _05278_ _05280_ _05284_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nand3_1
X_12041_ _04822_ _05209_ _04808_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12874_ _06109_ net277 _06100_ _06107_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__or4_4
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _04971_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__and2_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _04896_ _04897_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _03138_ _03153_ _03151_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__a21oi_2
X_11687_ _04817_ _04819_ _04820_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10638_ _03048_ _03049_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10569_ _02968_ _03595_ _02970_ _02972_ _02967_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a32o_2
X_12308_ _05160_ _05501_ _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12239_ _05073_ _05072_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07780_ _00680_ _00681_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__nor2_1
X_06800_ _06112_ _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__nor2_1
Xinput4 data_in[102] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_06731_ net105 VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09450_ _02365_ _02366_ _02302_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08401_ _01299_ _01300_ _01291_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__a21o_1
X_06662_ _04084_ _04095_ _04611_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__a21o_1
X_06593_ _03853_ _02492_ _03864_ _02503_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a22o_1
X_09381_ _01038_ _01620_ _01621_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08332_ _06284_ _06253_ _01230_ _01231_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__nand4_2
XFILLER_0_74_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08263_ _01142_ _00657_ _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07214_ _00114_ _00115_ net316 VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__a21oi_2
X_08194_ _01066_ _01067_ _01093_ _01094_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07145_ _00047_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07076_ net235 _05969_ _06001_ _03886_ _05980_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07978_ net52 net62 VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__and2_1
X_09717_ _02578_ _02659_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__nand3_2
X_06929_ net160 VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__clkbuf_4
X_09648_ _01981_ _02000_ _02001_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__nor3_2
XFILLER_0_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _02507_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__or2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _05810_ _05811_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__nor2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11610_ _00270_ _01754_ _04282_ _04279_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__a31oi_4
X_11541_ _01666_ _01652_ _03006_ _00550_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11472_ _04569_ _04585_ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10423_ _02818_ _02827_ _02826_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__a21o_1
X_10354_ _03355_ _03356_ _03357_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10285_ _02616_ _03281_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__nor2_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _04803_ _05190_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12857_ _06097_ _06094_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11808_ _04511_ _04954_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12788_ _05954_ _05965_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11739_ _04846_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08950_ _01817_ _01818_ _01848_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__o21ba_1
X_08881_ _06130_ _01777_ _01779_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__o2bb2a_1
X_07901_ _00419_ _00141_ _00581_ _00582_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__o211ai_4
X_07832_ _00660_ _00661_ _00733_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07763_ net136 VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__buf_2
X_09502_ _02422_ _02423_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__xnor2_1
X_06714_ net175 VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07694_ _06236_ _06240_ _00595_ _00596_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__o211ai_4
X_09433_ _01665_ _01669_ _01668_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__a21bo_1
X_06645_ net25 VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09364_ net229 net221 net222 net228 VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__a22o_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _00705_ _01215_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__xnor2_1
X_06576_ _03513_ _03678_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09295_ _01601_ _01691_ _01692_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08246_ _04227_ _00617_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__a21oi_1
X_08177_ _02789_ _03106_ _00550_ net212 VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__nand4_1
XFILLER_0_50_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07128_ _00029_ _00030_ _05246_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07059_ net6 net7 net254 net255 VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__nand4_2
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10070_ _02109_ _02379_ _02378_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10972_ _00956_ _00910_ net119 _00454_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12711_ _05803_ _05939_ _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__a21o_1
X_12642_ _05866_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12573_ _05781_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11524_ _00516_ _03580_ _04643_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11455_ _04115_ _04120_ _04114_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a21o_1
X_10406_ _03412_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__xnor2_2
X_11386_ _03986_ _04010_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10337_ _03336_ _03338_ _03339_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand3_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _01293_ net144 VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__and2_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _05150_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__xnor2_1
X_10199_ _02555_ _02556_ _02548_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09080_ _01363_ _01372_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__or2_1
X_08100_ net187 VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__buf_2
Xinput40 data_in[135] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
X_08031_ _00930_ _00931_ _00919_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput73 data_in[165] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
Xinput51 data_in[145] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput62 data_in[155] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput95 data_in[185] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 data_in[175] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09982_ _01023_ _02950_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08933_ _01829_ _01832_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08864_ _01729_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__xnor2_2
X_07815_ net96 net88 net90 net95 VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08795_ _01693_ _01694_ _01101_ net323 VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__a211o_1
X_07746_ _00645_ _00646_ _02207_ _00647_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09416_ _03095_ net1 net56 net67 VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__nand4_2
XFILLER_0_66_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07677_ _00577_ _00578_ _00135_ net297 VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06628_ _04227_ _02317_ _04238_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__and3_1
X_09347_ _02250_ _02252_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nand3_2
X_06559_ _03326_ _03491_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09278_ _01559_ _02177_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__nand3_1
XFILLER_0_132_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08229_ _01129_ _01130_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11240_ _04330_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__xnor2_2
X_11171_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10122_ _03093_ _03094_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__a21oi_1
X_10053_ _02337_ _02357_ _02356_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10955_ _03918_ _04017_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nand2_1
X_10886_ _03347_ _03350_ _03349_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12625_ _05817_ _05818_ _05848_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__nor3_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ _05543_ _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11507_ _03574_ _04124_ _04122_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12487_ _05689_ _05381_ _05698_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__nand3_1
XFILLER_0_110_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11438_ _00454_ _02132_ _04548_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11369_ _04459_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08580_ _00423_ _01480_ _00944_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__o21ai_1
X_07600_ _00072_ _00501_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07531_ _05498_ _05520_ _00432_ _00433_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07462_ _06380_ _00364_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07393_ _00293_ _00294_ _00295_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__or3_2
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09201_ _02056_ _02057_ _02099_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09132_ _02028_ _02031_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09063_ _01899_ _01961_ _01962_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__or3_4
XFILLER_0_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08014_ _00914_ _00915_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09965_ net193 net188 VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08916_ _01234_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__xor2_1
X_09896_ _03381_ net181 _02164_ _03546_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a22oi_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _01744_ _01746_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__xor2_1
X_08778_ _01675_ _01676_ _01677_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07729_ _00264_ _00287_ _00629_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__nor3_1
X_10740_ _00200_ net101 VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10671_ _02466_ _03100_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12410_ _05613_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12341_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12272_ _04974_ _05108_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__a21o_1
X_11223_ _03774_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__xor2_1
X_11154_ _03076_ _03077_ _03680_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21o_1
X_11085_ _04140_ _04160_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__and2_1
X_10105_ _03083_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nand2_2
Xinput252 data_in[96] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xinput241 data_in[86] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_2
Xinput230 data_in[76] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
X_10036_ _03003_ _03010_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ _04737_ _04755_ _04753_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10938_ _00431_ _01443_ _02064_ _06424_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_58_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10869_ _03340_ _03341_ _03344_ _02697_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a31o_2
XFILLER_0_39_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12608_ _05825_ _05830_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12539_ _05539_ _05561_ _05559_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09750_ _03864_ net246 net241 net242 VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__and4_1
X_06962_ _04314_ net124 net125 _02218_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09681_ _02612_ _02620_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__xnor2_1
X_08701_ _01033_ _01043_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__and2_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08632_ _00982_ _01531_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__nand3_1
X_06893_ _04270_ _04556_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__nand2_1
X_08563_ _01429_ _01463_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__xor2_2
X_08494_ _01384_ _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__xnor2_2
X_07514_ _06402_ _00414_ _00415_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__nor3_1
X_07445_ _06364_ _00347_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07376_ _00269_ _00276_ _00277_ _00278_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09115_ _02012_ _02013_ _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09046_ _06311_ _01293_ _01943_ _01944_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__and4_2
XFILLER_0_103_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09948_ _02908_ _02909_ _02913_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__o211ai_2
X_09879_ _02836_ _02837_ _02831_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__a21o_1
X_11910_ _01653_ _01629_ _02329_ _01051_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a22oi_1
X_12890_ clknet_1_0__leaf_clk _00014_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dfxtp_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11841_ _04549_ _04551_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__nand2_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _04461_ _04463_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _03748_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__xnor2_2
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10654_ _03687_ _03688_ _00166_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10585_ _03611_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12324_ _05274_ _05348_ _05519_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12255_ _05080_ _05083_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__nand2_1
X_11206_ _03917_ _04020_ _04019_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__a21o_2
X_12186_ _04612_ _05039_ _05037_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__a21bo_1
X_11137_ _04022_ _04219_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__xnor2_4
X_11068_ _00080_ _04123_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__nand2_1
X_10019_ _02312_ _02314_ _02313_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07230_ _00131_ _00132_ _00095_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o21ai_1
X_07161_ _02745_ _00062_ _00063_ _00064_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07092_ _06112_ _06404_ _06405_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__nand3_2
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09802_ _02084_ _02086_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__nand2_1
X_07994_ _00869_ _00895_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__xnor2_1
X_09733_ _02674_ _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__xor2_1
X_06945_ _06257_ _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__nor2_1
X_09664_ _02599_ _02600_ _02595_ _01946_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a211o_1
X_06876_ _06189_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__and2_1
X_09595_ _06253_ _00672_ _02524_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__a22o_1
X_08615_ _01482_ _01483_ _01513_ _01514_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _01445_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08477_ _01376_ _01377_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07428_ _00329_ _00330_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__or2_2
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07359_ _00261_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10370_ _02725_ _02738_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09029_ _01321_ _01329_ _01328_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ _05207_ _05208_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12873_ _06109_ _06100_ _06107_ net277 VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__o31ai_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04891_ _04970_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__or2_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _02694_ _01367_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _03200_ _03201_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__o21a_2
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11686_ _00665_ _01872_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10637_ _03316_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10568_ _02969_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10499_ _03517_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nor2_2
X_12307_ _01157_ _01754_ _05159_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__and3_1
X_12238_ _05406_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__xor2_4
X_12169_ _05028_ _05051_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
Xinput5 data_in[103] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06730_ _03568_ _03634_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__or2_1
X_06661_ _04084_ _04095_ _04611_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__nand3_2
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08400_ _01291_ _01299_ _01300_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__nand3_2
X_06592_ net244 VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__clkbuf_4
X_09380_ _02288_ _02289_ _01619_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08331_ _06284_ net97 _01230_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08262_ _01161_ _01162_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__nand2_1
X_07213_ _00114_ _00115_ _00116_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08193_ _01066_ _01067_ _01093_ _01094_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__nor4_1
XFILLER_0_104_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07144_ _03348_ net184 _00047_ net191 VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07075_ _06387_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07977_ net55 VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_4
X_09716_ _02656_ _02658_ _01961_ _02579_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__a211o_1
X_06928_ _06195_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06859_ _03941_ _04106_ _06173_ _02459_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__a22oi_1
X_09647_ _01934_ _01955_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09578_ _02505_ _02506_ _01837_ _01839_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__a211oi_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _00891_ _00893_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__nand2_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11540_ _04182_ _04185_ _04184_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11471_ _04583_ _04584_ _04570_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10422_ _02806_ _02808_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nand2_1
X_10353_ _03355_ _03356_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10284_ _02616_ _03281_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12023_ _04781_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12856_ net273 VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__inv_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _01487_ _02064_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__and3_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12787_ _05953_ _05951_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11738_ _04848_ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11669_ _04800_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08880_ net165 net166 net163 net164 VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07900_ _00799_ _00800_ _00638_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__o21a_1
X_07831_ _00692_ _00732_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__xnor2_2
X_07762_ _00207_ _00218_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__or2_1
X_09501_ _06243_ net171 VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06713_ net100 VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07693_ _00593_ _00594_ _00169_ _00154_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__a211o_1
X_09432_ _02345_ _02346_ _02344_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__a21o_1
X_06644_ net16 VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__buf_2
X_09363_ _02270_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06575_ _03656_ _03667_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ _01213_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09294_ _02194_ _02195_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08245_ _01144_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__nor2_1
X_08176_ net12 net190 VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07127_ _05246_ _00029_ _00030_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07058_ _06369_ _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10971_ _04026_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__xor2_4
XFILLER_0_97_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12710_ _05940_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12641_ _05686_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12572_ _05790_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__nor2_2
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11523_ _00086_ _01617_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11454_ _04076_ _04078_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10405_ _02771_ _03413_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11385_ _03987_ _04009_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10336_ _03336_ _03338_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a21o_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _06171_ _06319_ net146 net147 VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__nand4_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _05151_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__xnor2_4
X_10198_ _02522_ _02530_ _02529_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12839_ _06079_ _06080_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 data_in[126] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08030_ _00919_ _00930_ _00931_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput41 data_in[136] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xinput63 data_in[156] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput52 data_in[146] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput85 data_in[176] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xinput74 data_in[166] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xinput96 data_in[186] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
X_09981_ net220 net231 net232 net219 VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _01830_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08863_ _01730_ _01762_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07814_ _00231_ _00232_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08794_ _01101_ net294 _01693_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o211a_1
X_07745_ net29 VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__buf_2
X_09415_ _03095_ net56 net67 net1 VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__a22o_1
X_07676_ _00135_ net297 _00577_ _00578_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06627_ _04227_ _02317_ _04238_ _02328_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09346_ _01582_ _01592_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__a21o_1
X_06558_ _03469_ _03480_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09277_ _02175_ _02176_ _02168_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__a21o_1
X_06489_ net167 VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08228_ _00606_ _00607_ _00605_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08159_ _01058_ _01059_ _01060_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11170_ _03738_ _03697_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10121_ _03101_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__xor2_1
X_10052_ _03013_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10954_ _03918_ _04017_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nor2_1
X_10885_ _03940_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__or2_2
X_12624_ _05817_ _05818_ _05848_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12555_ _04775_ _05524_ _05525_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11506_ _04623_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12486_ _05689_ _05381_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11437_ _00956_ _00910_ _01520_ _01484_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__nand4_2
X_11368_ _04471_ _04472_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10319_ _02704_ _02719_ _02718_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__a21bo_2
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11299_ _04394_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__xnor2_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07530_ _02657_ _03590_ _06424_ _00431_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__nand4_1
XFILLER_0_88_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07461_ _00361_ _00363_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07392_ _06312_ _00292_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__and2b_1
X_09200_ _02097_ _02098_ _02059_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09131_ _02029_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09062_ _01959_ _01960_ _01900_ _01427_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08013_ net79 _06424_ _00912_ _00913_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__nand4_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09964_ net192 net189 VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__nand2_1
X_08915_ _01806_ _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__xnor2_1
X_09895_ _02202_ _02209_ _02208_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__a21o_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _01143_ _01147_ _01148_ _01745_ _01151_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__o32a_1
X_08777_ _01675_ _01676_ _01677_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07728_ _00264_ _00287_ _00629_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07659_ _00558_ _00559_ _00560_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _03157_ _03131_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09329_ _01589_ _01590_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12340_ _05192_ _05195_ _05536_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12271_ _05105_ _05107_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11222_ _04310_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ _03061_ _03683_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__and2_1
Xinput220 data_in[67] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_4
X_11084_ _04140_ _04160_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nor2_1
X_10104_ _02445_ _02417_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__or2b_1
Xinput242 data_in[87] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
Xinput253 data_in[97] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput231 data_in[77] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_4
X_10035_ _03003_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _04764_ _04888_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10937_ _03409_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10868_ _02676_ _03330_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a21o_2
X_12607_ _05825_ _05830_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10799_ _03768_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__xor2_4
XFILLER_0_53_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12538_ _05497_ _05506_ _05504_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12469_ _05385_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06961_ _02218_ _04314_ _06152_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nand4_1
X_09680_ _02618_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__and2b_1
X_08700_ _01599_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__nand2_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08631_ _01529_ _01530_ _01523_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__a21o_1
X_06892_ _02415_ _04600_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08562_ _01460_ _01462_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08493_ _01392_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07513_ _00414_ _00415_ _06402_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__o21a_1
X_07444_ _00345_ _00346_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07375_ _00274_ _00275_ _06267_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__or3b_2
X_09114_ _01387_ _01389_ _01388_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09045_ _06311_ _01293_ _01943_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_115_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09947_ _00049_ _01567_ _02911_ _02912_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__nand4_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09878_ _02831_ _02836_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__nand3_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _01140_ _01167_ _01169_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__a21o_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _04988_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__xnor2_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _04912_ _04913_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _03750_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__xnor2_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ _03068_ _03071_ _03067_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10584_ _02988_ _02990_ _02989_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12323_ _05347_ _05276_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12254_ _04639_ _05044_ _05043_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11205_ _03848_ _03912_ _03910_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__a21o_2
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12185_ _05013_ _05014_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__nor2_1
X_11136_ _04215_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__xor2_4
X_11067_ _04141_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__or2_1
X_10018_ _02988_ _02989_ _02990_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11969_ _04253_ _04718_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07160_ _03381_ _03392_ _05191_ _05202_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__nand4_4
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07091_ _06402_ _06403_ _05619_ _05663_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09801_ _02113_ _02124_ _02123_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09732_ _02675_ _02676_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__or2_1
X_07993_ _00893_ _00894_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__nand2_1
X_06944_ _02251_ _06253_ _06255_ _06256_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09663_ _02595_ _01946_ _02599_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_97_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06875_ _06170_ _03974_ _06188_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09594_ _04413_ _06254_ net92 _01858_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__nand4_2
X_08614_ _01482_ _01483_ _01513_ _01514_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__nand4_4
X_08545_ net68 net59 _01443_ _01444_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08476_ _01360_ _01375_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07427_ _06396_ _06399_ _00327_ _00328_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07358_ _00259_ _00260_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ _00170_ _00191_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__xnor2_1
X_09028_ _01925_ _01926_ _01917_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12872_ net320 _06108_ _06110_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11823_ _04891_ _04970_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__nand2_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _01385_ _01987_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11685_ _00677_ _01264_ _01250_ _03210_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__and4_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _03187_ _03202_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10636_ _03666_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__xor2_4
XFILLER_0_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10567_ _02969_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10498_ _03515_ _03516_ _03432_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _02464_ _01754_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12237_ _05424_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand2_2
X_12168_ _05001_ _05021_ _05019_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a21o_1
X_11119_ _03629_ _03643_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a21o_1
X_12099_ _04937_ _04968_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__a21bo_1
Xinput6 data_in[104] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_06660_ _02415_ _04600_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06591_ net236 VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__clkbuf_4
X_08330_ _04413_ _06254_ net90 net91 VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nand4_2
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08261_ _01159_ _01160_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07212_ net1 net12 _04950_ _03128_ _04939_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08192_ _01091_ _01092_ _00561_ _00563_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07143_ net185 VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07074_ _03853_ _05969_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07976_ _00876_ _00877_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__nor2_1
X_09715_ _01961_ net293 _02656_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__o211ai_4
X_06927_ _06239_ _06240_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__nor2_1
X_09646_ _02003_ _02054_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06858_ _06172_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06789_ _02503_ _05969_ _05991_ _06001_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_93_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09577_ _01837_ _01839_ _02505_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o211a_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _01427_ _01428_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__and2_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _01359_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11470_ _04570_ _04583_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10421_ _02891_ _02942_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10352_ _02705_ _02713_ _02711_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10283_ _03279_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__xor2_1
X_12022_ _05187_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__xnor2_2
X_12855_ _06096_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__clkbuf_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _01488_ _01443_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__and2_1
X_12786_ _06018_ _06025_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__xor2_1
X_11737_ _04850_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__xor2_2
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11668_ _00672_ _03180_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10619_ _03002_ _03032_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11599_ _04723_ _04724_ _04725_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07830_ _00730_ _00731_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__nor2_1
X_07761_ _00208_ _00217_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__or2_1
X_06712_ _05158_ _05169_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__or2_1
X_09500_ _02420_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__nand2_1
X_07692_ _00169_ _00154_ _00593_ _00594_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__o211ai_4
X_09431_ _02344_ _02345_ _02346_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__nand3_1
X_06643_ _04413_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09362_ net217 net233 VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06574_ _02701_ _03645_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08313_ _01211_ _01212_ net85 net101 VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09293_ _02192_ _02193_ _02111_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08244_ net159 net160 net169 net170 VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__and4_1
X_08175_ _01073_ _01076_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07126_ _02635_ _03546_ _05389_ _06437_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__and4_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07057_ _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07959_ _00844_ _00860_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__xnor2_1
X_10970_ _04027_ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__xor2_4
X_09629_ _02562_ _02563_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12640_ _01488_ _01443_ _02799_ _02064_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__and4_2
XFILLER_0_38_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12571_ _05789_ _05784_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__and2b_1
X_11522_ _04640_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11453_ _04060_ _04078_ _04079_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10404_ _02774_ _02775_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11384_ _04455_ _04489_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10335_ net239 net249 VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__and2_1
X_10266_ net151 net146 net147 net150 VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a22o_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12005_ _05152_ _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10197_ _03170_ _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12838_ _06079_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__nand2_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _05916_ _05926_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput31 data_in[127] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
Xinput20 data_in[117] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_4
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 data_in[157] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
Xinput42 data_in[137] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput53 data_in[147] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput86 data_in[177] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xinput97 data_in[187] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
Xinput75 data_in[167] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09980_ net219 net220 net232 VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__and3_1
X_08931_ net85 net102 net22 net24 VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08862_ _01731_ _01761_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__xnor2_4
X_07813_ _00702_ _00713_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__and2_1
X_08793_ _01691_ _01692_ _01601_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_74_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07744_ _00644_ net160 net168 _00642_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07675_ _00575_ _00576_ _00504_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__a21o_1
X_09414_ net40 VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06626_ net166 VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09345_ _01591_ _01583_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__and2b_1
X_06557_ _02767_ _03458_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06488_ net182 VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__clkbuf_4
X_09276_ _02168_ _02175_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__nand3_2
XFILLER_0_35_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08227_ net281 _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08158_ _03084_ _00097_ _00534_ _00533_ _00107_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07109_ net76 net77 net70 net71 VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__and4_1
X_08089_ net183 net184 _00989_ _00480_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__nand4_1
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10120_ _02422_ _02423_ _02421_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o21ai_1
X_10051_ _03026_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__xor2_4
XFILLER_0_100_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10953_ _03980_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__xnor2_1
X_10884_ _03938_ _00830_ _01385_ _03937_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__and4b_1
XFILLER_0_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ _05836_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xnor2_1
X_12554_ _05544_ _05545_ _05207_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11505_ _04619_ _04620_ _04621_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12485_ _05690_ _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11436_ _00910_ _01520_ _01484_ _00956_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__a22o_1
X_11367_ _04467_ _04469_ _04470_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10318_ _02671_ _02681_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__a21bo_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11298_ _01293_ _02615_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and3_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10249_ _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07460_ _06372_ _06374_ _06376_ _00362_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07391_ _04139_ _06311_ _00291_ _02383_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09130_ _01396_ _01398_ _01399_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09061_ _01900_ _01427_ _01959_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08012_ _05520_ _06424_ _00912_ _00913_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09963_ _02268_ _02271_ _02269_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08914_ _01807_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09894_ _02175_ _02177_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _01150_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__inv_2
X_08776_ _01077_ _01085_ _01084_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07727_ _00627_ _00628_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__and2_1
X_07658_ _00558_ _00559_ _00560_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__nand3_4
XFILLER_0_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07589_ _05115_ _05093_ _00490_ _00491_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06609_ _04029_ _04040_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and2_1
X_09328_ _02231_ _02232_ _02211_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09259_ _01533_ _01536_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12270_ _05349_ _05461_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11221_ _04307_ _04308_ _04309_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__o21bai_1
X_11152_ _04233_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__xor2_2
XFILLER_0_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10103_ _02444_ _02418_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__or2b_1
Xinput210 data_in[58] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlymetal6s2s_1
X_11083_ _04152_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__xnor2_1
Xinput254 data_in[98] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_4
Xinput221 data_in[68] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_4
Xinput232 data_in[78] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_2
Xinput243 data_in[88] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__buf_2
X_10034_ _03004_ _03008_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11985_ _04765_ _04887_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__and2_1
X_10936_ net71 net72 net83 net84 VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__and4_1
X_10867_ _03325_ _03329_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12606_ _05828_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _03845_ _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12537_ _05521_ _05581_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12468_ _05676_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11419_ _04438_ _04527_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12399_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06960_ net125 VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__buf_2
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06891_ _06203_ _06204_ _04084_ _04622_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__o211a_1
X_08630_ _01523_ _01529_ _01530_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08561_ _00403_ _00896_ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08492_ _01390_ _01391_ _01386_ _00837_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07512_ net296 _00413_ _00341_ _00042_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__o211a_1
X_07443_ _00342_ _06392_ _00344_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09113_ _02009_ _02010_ _02011_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__nand3_1
X_07374_ _06267_ net308 _00276_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09044_ _06171_ net151 net143 _00774_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__nand4_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ _00047_ _01567_ _02911_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09877_ _02832_ _02834_ _02835_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__nand3_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _01708_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__inv_2
X_08759_ _03095_ _01072_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__nand2_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _00850_ _02019_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__nand2_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _03751_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10652_ _03685_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__nor2_1
X_10583_ _03609_ _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12322_ _05265_ _05267_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12253_ _05441_ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__or2_2
X_11204_ _04258_ _04291_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12184_ _05365_ _05366_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__and2_2
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11135_ _03519_ _03661_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a21oi_2
X_11066_ net221 net222 net231 net232 VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__and4_1
X_10017_ _02988_ _02989_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11968_ _04236_ _04719_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__and2_1
X_10919_ _03936_ _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__xor2_2
X_11899_ _01072_ _03019_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__nand2_2
XFILLER_0_128_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07090_ _05619_ _05663_ _06402_ _06403_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09800_ _02079_ _02091_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__or2_2
X_07992_ _00891_ _00892_ _00870_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__a21o_1
X_09731_ net236 net237 net250 net251 VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__and4_2
X_06943_ net85 _06253_ _06255_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09662_ _02596_ _02597_ _02598_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__nand3_1
X_06874_ _06170_ _03974_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__o21ai_2
X_09593_ _06254_ net92 _01858_ _04413_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__a22o_1
X_08613_ _01510_ _01511_ _01512_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08544_ net68 _01443_ _01444_ net59 VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__a22oi_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08475_ _01360_ _01375_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07426_ _00327_ _00328_ _06396_ _06399_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07357_ _00237_ _00258_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09027_ _01917_ _01925_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07288_ _00189_ _00190_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09929_ net175 net145 net156 net174 VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12871_ _06109_ _06100_ _06107_ _02185_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__o31a_1
X_11822_ _04892_ _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _04459_ _04472_ _04471_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11684_ _01264_ _01250_ _03210_ _00677_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__a22oi_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10704_ _03135_ _03155_ _03742_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_126_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10635_ _02793_ _03047_ _03668_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10566_ _03591_ _03592_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__xnor2_4
X_12305_ _05198_ _05183_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10497_ _03432_ _03515_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__and3_1
X_12236_ _05408_ _05409_ _05423_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__or3_1
X_12167_ _05274_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__xor2_1
X_11118_ _03642_ _03640_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__and2b_1
X_12098_ _04965_ _04967_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nand2_1
Xinput7 data_in[105] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11049_ net233 VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06590_ _02481_ _03787_ _03809_ _03831_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__a22o_2
XFILLER_0_47_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08260_ _01159_ _01160_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__nand2_2
X_07211_ _00112_ _00113_ _00111_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__a21o_1
X_08191_ _00561_ _00563_ net306 _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07142_ _00045_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07073_ _06384_ _06385_ _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07975_ _00871_ _00875_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__nor2_1
X_09714_ _02654_ _02655_ _02581_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__a21o_1
X_06926_ _06208_ _06238_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__nor2_2
X_06857_ net210 VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__buf_2
X_09645_ _02053_ _02052_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06788_ net235 _05969_ _05991_ _06001_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09576_ _06159_ _01835_ _02502_ _02504_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__nand4_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _01425_ _01426_ _01378_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08458_ _00809_ _00811_ _00812_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07409_ _00310_ _00309_ _00296_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_108_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08389_ _04128_ net139 _00749_ _01288_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10420_ _02882_ _02884_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10351_ _03353_ _03354_ _03346_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10282_ _06086_ net216 VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nand2_1
X_12021_ _04776_ _04779_ _04777_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__o21ba_1
X_12854_ _02174_ _06093_ _06094_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _04949_ _04951_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__xnor2_4
X_12785_ _06019_ _06024_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__xnor2_1
X_11736_ _04864_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__xor2_4
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ _04798_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10618_ _03029_ _03030_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__and2_1
X_11598_ _04723_ _04724_ _00166_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10549_ net220 net221 net231 net232 VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12219_ _05403_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__xnor2_4
X_07760_ _06323_ _00219_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06711_ _05137_ _05147_ _05082_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__a21oi_1
X_09430_ _03106_ net223 net234 _02789_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__a22o_1
X_07691_ _00591_ _00592_ _00192_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__a21o_1
X_06642_ net95 VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09361_ _02268_ _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06573_ _02701_ _03645_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08312_ net85 net101 _01211_ _01212_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o2bb2a_1
X_09292_ _02111_ _02192_ _02193_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__nand3_1
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08243_ net160 net169 _00171_ net159 VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08174_ _01074_ _01075_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07125_ _00028_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__inv_2
X_07056_ net253 net252 net8 net9 VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ _00858_ _00859_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__xnor2_1
X_07889_ _00788_ _00789_ _00381_ _00738_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__o211a_1
X_06909_ _06223_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
X_09628_ net132 net128 VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09559_ net27 net20 net21 net26 VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a22o_1
X_12570_ _05784_ _05789_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__and2b_2
XFILLER_0_93_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11521_ _00507_ _04123_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11452_ _04547_ _04564_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10403_ _02774_ _02775_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__nor2_1
X_11383_ _04486_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__xnor2_2
X_10334_ net247 net248 net240 net241 VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nand4_1
X_10265_ _03259_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__xor2_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ _03184_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__nor2_1
X_12004_ _05154_ _05168_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12837_ _06071_ _06074_ _06069_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12768_ _05938_ _05946_ _05944_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__o21a_1
X_11719_ _00774_ _02592_ _04855_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12699_ _05852_ _05881_ _05850_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__a21oi_2
Xinput21 data_in[118] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xinput10 data_in[108] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput54 data_in[148] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xinput43 data_in[138] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xinput32 data_in[128] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput76 data_in[168] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput87 data_in[178] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
Xinput98 data_in[188] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xinput65 data_in[158] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
XFILLER_0_40_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08930_ net85 net24 net102 net22 VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nand4_1
X_08861_ _01733_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__xnor2_4
X_07812_ _00702_ _00713_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08792_ _01601_ _01691_ _01692_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07743_ net168 net160 _00643_ _00644_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07674_ _00504_ _00575_ _00576_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__nand3_4
X_09413_ _03095_ _01072_ _01662_ _01661_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a31o_1
X_06625_ net158 VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09344_ _02248_ _02249_ _02235_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06556_ _02767_ _03458_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06487_ net191 VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__clkbuf_4
X_09275_ _02172_ _02173_ _02169_ _01528_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08226_ _00611_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__xnor2_1
X_08157_ _01056_ _01057_ _01055_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07108_ _06419_ _06420_ _05455_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__o21a_1
X_08088_ net184 _00989_ _00480_ net183 VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07039_ _05783_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10050_ _02343_ _02352_ _02351_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_98_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10952_ _04013_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10883_ _01385_ _00830_ _03937_ _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_78_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12622_ _05837_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12553_ _05523_ _05528_ _05532_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11504_ _04619_ _04620_ _04621_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ _05694_ _05695_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11435_ _04544_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__nor2_2
X_11366_ _04467_ _04469_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11297_ _06319_ _01309_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__nand2_1
X_10317_ _02680_ _02672_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__or2b_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10248_ _03203_ _03241_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nor2_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ _02500_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07390_ _00292_ _06312_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09060_ _01957_ _01958_ _01901_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08011_ _02657_ _03590_ _00431_ net73 VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__nand4_4
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09962_ _02241_ _02243_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08913_ _01253_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__xnor2_1
X_09893_ _01559_ _02177_ _02178_ _02181_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__a31o_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _01742_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__xnor2_1
X_08775_ _01673_ _01674_ _01664_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07726_ _00281_ _00284_ _00626_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__or3_1
X_07657_ _00110_ _00118_ net315 VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__o21bai_2
X_07588_ net191 net192 _00047_ _00489_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06608_ _02602_ _04018_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06539_ _03249_ _03271_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09327_ _02211_ _02231_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__nor3_1
XFILLER_0_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ _02155_ _02156_ _02126_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09189_ _02087_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__or2b_1
X_08209_ _00905_ _00906_ _01109_ _01110_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__nor4_1
XFILLER_0_114_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11220_ _04307_ _04308_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__or3b_2
XFILLER_0_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ _03079_ _03679_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10102_ _02453_ _02664_ _02663_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__a21o_2
Xinput200 data_in[49] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
Xinput211 data_in[59] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
X_11082_ _04156_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__xor2_1
Xinput244 data_in[89] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_4
Xinput233 data_in[79] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_2
Xinput222 data_in[69] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
X_10033_ _03005_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand2_1
Xinput255 data_in[99] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_2
X_11984_ _04734_ _04758_ _04760_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10935_ _06347_ _02765_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10866_ _03345_ _03360_ _03358_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a21o_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _05656_ _05826_ _05668_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__nor3_1
XFILLER_0_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10797_ _03769_ _03242_ _03844_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nor3_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12536_ _05582_ _05518_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12467_ _05430_ _05452_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_81_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11418_ _04438_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12398_ _05598_ _05600_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11349_ _03328_ _03931_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06890_ _04084_ _04622_ _06203_ _06204_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08560_ _00869_ _00893_ _00894_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__and3_1
X_08491_ _01386_ _00837_ _01390_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__o211ai_1
X_07511_ _00341_ _00042_ net296 _00413_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_119_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07442_ _00342_ _06392_ _00344_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07373_ _00274_ _00275_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__or2_1
X_09112_ _02009_ _02010_ _02011_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09043_ net151 net143 net144 net150 VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09945_ _00989_ net186 _00480_ net187 VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__nand4_1
X_09876_ _02832_ _02834_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__a21o_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _01139_ _01169_ _01170_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o31ai_4
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _01657_ _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__nor2_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08689_ _01004_ _01006_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07709_ _00603_ _00600_ _00599_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__a21oi_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10720_ _03759_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__nand2_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10651_ net285 _03684_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10582_ _04862_ net44 net39 net40 VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12321_ _05233_ _05269_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12252_ _05032_ _05440_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11203_ _04261_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__xnor2_2
X_12183_ _05354_ _05364_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nand2_1
X_11134_ _03658_ _03660_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nor2_1
X_11065_ net222 net231 _01603_ net221 VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__a22oi_1
X_10016_ net44 net38 VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11967_ _05128_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10918_ _03976_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11898_ _04661_ _04668_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__and2_2
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10849_ _03857_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12519_ net263 _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07991_ _00870_ _00891_ _00892_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__nand3_1
X_09730_ _05980_ _01367_ _01987_ _03853_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__a22oi_1
X_06942_ _04413_ net87 _06254_ net86 VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09661_ _02596_ _02597_ _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a21o_1
X_06873_ _06186_ _06187_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__nor2_2
X_09592_ _01855_ _01859_ _01856_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08612_ _01510_ _01511_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__nand3_4
X_08543_ net57 VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08474_ _00842_ _01374_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07425_ _00289_ _06326_ _00326_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__nand3_2
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07356_ _00237_ _00258_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07287_ _06337_ _06339_ _00188_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09026_ _01923_ _01924_ _01918_ _01919_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09928_ _02212_ _02216_ _02213_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__o21bai_1
X_09859_ _03590_ net79 _01488_ net75 VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12870_ net276 VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__inv_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _04937_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__xnor2_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04448_ _04449_ _04452_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11683_ _00201_ _01264_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__and2_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10703_ _03154_ _03136_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__and2b_1
X_10634_ _03045_ _03046_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10565_ _04906_ net49 VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nand2_2
X_12304_ _05197_ _05184_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10496_ _03512_ _03514_ _03433_ _02945_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12235_ _05408_ _05409_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12166_ _05276_ _05347_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__xnor2_1
X_11117_ _04190_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__xnor2_4
X_12097_ _05179_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__xor2_2
Xinput8 data_in[106] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
X_11048_ _03577_ _03587_ _03586_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07210_ _00111_ _00112_ _00113_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__nand3_1
X_08190_ _01089_ _01090_ _01071_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__o21a_1
X_07141_ _05180_ _05268_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07072_ net244 net237 net238 net243 VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07974_ _00871_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__and2_1
X_09713_ _02581_ _02654_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__nand3_2
X_06925_ _06208_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__and2_1
X_06856_ net150 VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__clkbuf_4
X_09644_ _01957_ _01959_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06787_ _03853_ _03864_ _05980_ _02492_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__a22o_1
X_09575_ _06159_ _01835_ _02502_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__a22o_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _01378_ _01425_ _01426_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__or3_2
XFILLER_0_65_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08457_ _00969_ _00971_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__or2_2
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07408_ _00296_ _00309_ _00310_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08388_ _04128_ _00749_ _01288_ _02394_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07339_ _02251_ _00238_ _00240_ _00241_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10350_ _03346_ _03353_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09009_ _01906_ _01907_ _01903_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10281_ _06086_ net215 _02623_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12020_ _02498_ _01784_ _04775_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a31o_1
X_12853_ _06092_ _06090_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__or2_1
X_11804_ _00879_ _01434_ _04502_ _04500_ _02765_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a32o_2
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12784_ _06020_ _06022_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__xor2_1
X_11735_ _04872_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__xor2_4
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _04794_ _04795_ _04797_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a21oi_1
X_10617_ _03619_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11597_ _04243_ _04247_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10548_ _00507_ net231 _01603_ _00080_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12218_ _05054_ _05062_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__a21oi_4
X_10479_ _03493_ _03494_ _03495_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12149_ _05327_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06710_ _05082_ _05137_ _05147_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__and3_1
X_07690_ _00192_ _00591_ _00592_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__nand3_2
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06641_ _04358_ _04369_ _02273_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a21o_1
X_09360_ net218 net219 net231 net232 VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06572_ _03568_ _03634_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__xor2_1
X_08311_ net86 net87 net98 net99 VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09291_ _02190_ _02191_ _02112_ _01599_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08242_ _00644_ _00646_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08173_ net179 net23 net34 net112 VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07124_ _03546_ _05389_ _06437_ _02635_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07055_ _03820_ _05882_ _06368_ net252 VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07957_ _00354_ _00360_ _00359_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__a21bo_1
X_06908_ _02185_ _06221_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__and3_1
X_07888_ _00381_ _00738_ _00788_ _00789_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09627_ net131 net129 VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__nand2_1
X_06839_ _04303_ _04314_ _06152_ _02218_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a22o_1
X_09558_ _01829_ _01831_ _01830_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__a21bo_1
X_08509_ net4 VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ _04638_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__nor2_1
X_09489_ _01733_ _01760_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11451_ _04561_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__xor2_4
X_11382_ _03960_ _03975_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__a21bo_1
X_10402_ _03407_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10333_ net248 net240 net241 net247 VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10264_ _06178_ net155 VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__nand2_1
X_10195_ _02507_ _03171_ _03182_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nor3_1
X_12003_ _05166_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12836_ net268 VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__inv_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12767_ _06003_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__nor2_1
X_11718_ _00749_ _01309_ _01288_ _02615_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nand4_2
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12698_ _05928_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput22 data_in[119] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
Xinput11 data_in[109] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_0_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11649_ _04778_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__xnor2_1
Xinput44 data_in[139] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput55 data_in[149] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput33 data_in[129] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput88 data_in[179] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
Xinput77 data_in[169] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 data_in[159] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_0_12_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput99 data_in[189] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
XFILLER_0_40_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_08860_ _01161_ _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__xnor2_4
X_07811_ _00243_ _00712_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__xnor2_1
X_08791_ net310 _01689_ _01690_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__a21oi_2
X_07742_ _02317_ net166 net161 net162 VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07673_ net299 _00574_ _00505_ _00133_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__o211ai_4
X_09412_ _01678_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06624_ _02536_ _04205_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09343_ _02235_ _02248_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__nand3_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06555_ _03436_ _03447_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09274_ _02169_ _01528_ _02172_ _02173_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__o211ai_2
X_06486_ _02635_ _02646_ _02657_ _02668_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08225_ _01125_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__nor2_1
X_08156_ _01055_ _01056_ _01057_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07107_ _05455_ _06419_ _06420_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__nor3_1
X_08087_ net194 VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07038_ _06344_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08989_ _01886_ _01887_ _01854_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10951_ _03387_ _03421_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10882_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ _05839_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12552_ _05589_ _05639_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__a21bo_1
X_11503_ _04141_ _04144_ _04142_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12483_ _05438_ _05442_ _05693_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11434_ _04536_ _04543_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__and2_1
X_11365_ _03945_ _03953_ _03951_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11296_ _04392_ _04393_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__xnor2_1
X_10316_ _02795_ _02887_ _02886_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__a21o_1
X_10247_ _03203_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__and2_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ _03164_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12819_ _06058_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08010_ net77 net72 net73 net76 VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap300 net324 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_1
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09961_ _02272_ _02927_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__o21a_1
X_08912_ _01810_ _01811_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09892_ _02159_ _02183_ _02184_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__nand3_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _01145_ _01148_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__or2_1
X_08774_ _01664_ _01673_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07725_ _00281_ _00284_ _00626_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07656_ _00556_ _00557_ _00547_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07587_ _03348_ _00049_ _00489_ _02712_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__a22oi_1
X_06607_ _02602_ _04018_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__or2_1
X_06538_ _03227_ _02855_ _03260_ _02866_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a22o_1
X_09326_ _02227_ _02228_ _02230_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09257_ _02126_ _02155_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__nand3_2
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06469_ _02470_ _02481_ _02492_ _02503_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__a22o_1
X_08208_ net291 _01108_ net314 net309 VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09188_ _02085_ _02086_ _02082_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08139_ _00511_ _01035_ _01040_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__and3_1
X_11150_ _03675_ _03677_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nor2_1
X_10101_ _02414_ _02447_ _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput201 data_in[4] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
X_11081_ _02969_ _03593_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__a21oi_1
Xinput245 data_in[8] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_4
Xinput234 data_in[7] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
Xinput223 data_in[6] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
Xinput212 data_in[5] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
X_10032_ _03095_ _04939_ net56 _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nand4_1
Xinput256 data_in[9] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_6
X_11983_ _05123_ _04729_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__or2b_1
X_10934_ _03988_ _03995_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10865_ _03323_ _03332_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__a21o_2
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12604_ _05656_ _05826_ _05668_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o21a_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10796_ _03769_ _03242_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _05511_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12466_ _05429_ _05427_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12397_ _05598_ _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nand2_2
X_11417_ _04491_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11348_ _03926_ _03929_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11279_ _03811_ _03843_ _03840_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__o21a_1
X_07510_ _00383_ _00384_ _00411_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__o21a_1
X_08490_ _01387_ _01388_ _01389_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__nand3_1
X_07441_ _02448_ _00343_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07372_ _00273_ _06130_ _06127_ _00271_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__and4b_1
X_09111_ net246 net240 VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ _01940_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09944_ net186 net195 net187 _00989_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__a22o_1
X_09875_ net107 net117 VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__and2_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _01138_ _01172_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__or2b_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _01651_ _01656_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__nor2_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _01587_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__xnor2_1
X_07708_ _00610_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
X_07639_ _00540_ _00541_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__nand2_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10650_ net285 _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09309_ net183 net182 net197 net198 VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__and4_1
X_10581_ _00097_ _01653_ _02329_ _04862_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12320_ _05491_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12251_ _05032_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11202_ _04263_ _04289_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__xnor2_2
X_12182_ _05354_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or2_1
X_11133_ _04092_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__xnor2_4
X_11064_ _03602_ _03617_ _03616_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__a21oi_1
X_10015_ _03194_ _04862_ net39 net40 VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__nand4_2
XFILLER_0_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11966_ _05124_ _05127_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10917_ _03362_ _03379_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a21boi_2
X_11897_ _05026_ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10848_ _03878_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__xor2_2
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10779_ _03823_ _03824_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12518_ _05730_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__xor2_2
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12449_ _05656_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07990_ _00889_ _00890_ _00428_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06941_ net86 _04413_ net87 _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__nand4_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09660_ _00291_ _01293_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06872_ _02394_ _06171_ _06185_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__a21oi_1
X_08611_ _00919_ _00931_ _00930_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__a21bo_1
X_09591_ _04424_ _06134_ _00672_ _01251_ _01811_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__a41o_1
X_08542_ net83 VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08473_ _00811_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__xor2_1
X_07424_ _00289_ _06326_ _00326_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__a21o_2
XFILLER_0_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07355_ _00256_ _00257_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ _06337_ _06339_ _00188_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09025_ _01918_ _01919_ _01923_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09927_ _02204_ _02206_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__nand2_1
X_09858_ net79 _01488_ _02799_ _03590_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__a22oi_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _02724_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__xor2_4
X_08809_ _01173_ _01708_ _01709_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__and3_2
X_11820_ _04965_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__xor2_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _04532_ _04597_ _04596_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__a21oi_2
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _03317_ _03430_ _03428_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11682_ _00291_ _02592_ _04390_ _04389_ _01309_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__a32o_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10633_ _03431_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10564_ _02982_ _02985_ _02983_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12303_ _01188_ _01754_ _05163_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10495_ _03433_ _02945_ _03512_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_121_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12234_ _05420_ _05421_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12165_ _05318_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__xor2_1
X_11116_ _03624_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__xor2_4
X_12096_ _05181_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__xnor2_2
X_11047_ _04116_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__xnor2_4
Xinput9 data_in[107] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11949_ _04701_ _04703_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07140_ _04730_ _05060_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__or2b_1
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07071_ net243 net244 net237 VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09712_ _02652_ _02653_ _02582_ _02583_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__o211ai_4
X_07973_ _00873_ _00874_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__nor2_1
X_06924_ _06236_ _06237_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__or2_1
X_09643_ _01899_ _01961_ _01962_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__nor3_1
X_06855_ _02525_ _03919_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09574_ _06284_ _00200_ _00238_ _00703_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__nand4_1
X_08525_ _01379_ _00862_ _01424_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__nor3_1
X_06786_ _05980_ _03886_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08456_ _00899_ _00901_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__nand2_1
X_08387_ net154 VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__buf_2
X_07407_ _00308_ _00306_ _00307_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07338_ _02196_ _04446_ _06261_ _00239_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__nand4_2
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07269_ _04227_ _02328_ _06227_ _00171_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__nand4_1
X_09008_ _01903_ _01906_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10280_ _06361_ net204 net213 net214 VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__and4_1
XFILLER_0_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _06092_ _06090_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _04947_ _04948_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__or2_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12783_ _05933_ _05949_ _06021_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__a21bo_1
X_11734_ _04411_ _04412_ _04415_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__a21o_2
XFILLER_0_95_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11665_ _04794_ _04795_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__and3_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10616_ _03644_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__xor2_4
XFILLER_0_71_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11596_ _04721_ _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__nor2_1
X_10547_ _02980_ _03000_ _02999_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_52_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10478_ _03493_ _03494_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__nand3_1
XFILLER_0_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12217_ _05063_ _05070_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12148_ _01488_ _02064_ _04510_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__and3_1
X_12079_ _00757_ _03859_ _01986_ _02626_ _01365_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__o2111a_1
X_06640_ _04380_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06571_ _03601_ _03623_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__nand2_1
X_08310_ net87 net98 net99 net86 VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__a22oi_1
X_09290_ _02112_ _01599_ _02190_ _02191_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08241_ _00259_ _00655_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08172_ net112 net179 net23 net34 VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07123_ net106 VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07054_ net9 VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07956_ _00856_ _00857_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__or2b_1
X_06907_ _06219_ _06220_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__or2_1
X_07887_ _00786_ _00787_ _00740_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__a21oi_2
X_09626_ _01938_ _01941_ _01939_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__o21bai_2
X_06838_ _06152_ _04336_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__nand2_1
X_06769_ _02569_ _05750_ _05772_ _05794_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09557_ _01821_ _01823_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__nor2_1
X_08508_ _05914_ _00822_ _01406_ _01407_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nand4_1
XFILLER_0_65_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09488_ _01730_ _01762_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08439_ _01337_ _01338_ _01307_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11450_ _04046_ _04054_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a21boi_4
X_11381_ _03973_ _03971_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__or2b_1
X_10401_ _03408_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10332_ _03320_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10263_ _00749_ _03257_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a21bo_1
X_12002_ _05155_ _05156_ _05165_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__nand3_1
X_10194_ _02507_ _03171_ _03182_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _06078_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__clkbuf_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12766_ _05997_ _05928_ _06002_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__and3_1
X_11717_ _01309_ _01288_ _02615_ _00749_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__a22o_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12697_ _05915_ _05927_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__or2_1
Xinput12 data_in[10] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
X_11648_ _00706_ _01784_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 data_in[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 data_in[13] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 data_in[12] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
X_11579_ _04531_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__xnor2_4
Xinput89 data_in[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_4
Xinput78 data_in[16] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput67 data_in[15] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput56 data_in[14] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_0_122_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08790_ _01688_ _01689_ _01690_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__and3_2
X_07810_ _00710_ _00711_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__or2_1
X_07741_ _00642_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__inv_2
X_07672_ _00505_ _00133_ net299 _00574_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__a211o_4
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06623_ _04183_ _04194_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__and2_2
X_09411_ _02303_ _02324_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09342_ _02246_ _02247_ _02236_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__a21o_1
X_06554_ _03359_ _03370_ _03403_ _03425_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_118_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09273_ _03381_ _01524_ _02170_ _02171_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand4_2
XFILLER_0_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06485_ _02679_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08224_ _00595_ _00597_ _01123_ _01124_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__a211oi_1
X_08155_ _03194_ _04862_ net36 _00543_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__nand4_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07106_ _06417_ _06418_ _05411_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08086_ net182 net196 VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07037_ _06348_ _06350_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08988_ _01854_ _01886_ _01887_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nor3_2
X_07939_ _00832_ _00840_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10950_ _03388_ _03420_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__and2b_1
X_10881_ _06383_ _00366_ _02694_ net242 VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__and4_1
X_09609_ _02540_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__nor2_2
X_12620_ _05357_ _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12551_ _05640_ _05587_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__or2b_1
X_11502_ _04145_ _04151_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12482_ _05438_ _05442_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11433_ _04536_ _04543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11364_ _04464_ _04465_ _04466_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nand3_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11295_ _00291_ _02592_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10315_ _02749_ _02788_ _02787_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10246_ _03237_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__xor2_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10177_ _00250_ _00706_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12818_ _06014_ _06017_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12749_ _05984_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap301 _01095_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_1
XFILLER_0_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09960_ _01610_ _01611_ _02276_ _02277_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08911_ _06253_ _00200_ _01808_ _01809_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09891_ _02849_ _02850_ _02814_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a21oi_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _01736_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__xnor2_1
X_08773_ _01670_ _01671_ _01672_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__a21o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07724_ _00178_ _00625_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__xnor2_1
X_07655_ _00547_ _00556_ _00557_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__nand3_2
X_06606_ _03996_ _04007_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07586_ net186 VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06537_ net227 VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__buf_2
X_09325_ _02227_ _02228_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__and3_2
XFILLER_0_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06468_ net235 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ _02153_ _02154_ _01508_ _01510_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08207_ net314 net309 net291 _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09187_ _02082_ _02085_ _02086_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08138_ _01037_ _01039_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__nand2_1
X_08069_ _00908_ _00969_ _00970_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__nor3b_1
X_11080_ _04906_ _04154_ _03591_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__and3_1
X_10100_ _02446_ _02416_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__and2b_1
Xinput202 data_in[50] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
X_10031_ net67 VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput224 data_in[70] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_4
Xinput235 data_in[80] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_2
Xinput213 data_in[60] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
Xinput246 data_in[90] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
Xinput257 reset VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_4
X_11982_ _05120_ _05122_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__or2_1
X_10933_ _03993_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10864_ _03324_ _03331_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10795_ _03811_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__xor2_1
X_12603_ _05658_ _05650_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12534_ _05513_ _05495_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12465_ _05664_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_4
X_12396_ _02731_ _02019_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__and3_1
X_11416_ _04522_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11347_ _04448_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11278_ _04346_ _04373_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__xnor2_2
X_10229_ _03214_ _03215_ _03220_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_89_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07440_ net204 VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07371_ _06127_ _06130_ _00272_ _00273_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__o2bb2a_1
X_09110_ _02492_ _03864_ net241 net242 VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__nand4_1
XFILLER_0_17_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09041_ net139 net155 VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09943_ net184 net196 _02221_ _02222_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__and4_1
X_09874_ net115 net116 net108 net109 VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__nand4_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _00166_ _01725_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__nor2_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _01651_ _01656_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__and2_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ net193 _00489_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nand2_1
X_07707_ _02185_ _00608_ _00609_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__and3_1
X_07638_ _00103_ _00539_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__or2_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ _05191_ _05202_ _00059_ _03392_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09308_ net183 net197 net198 net182 VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10580_ _03606_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09239_ _02137_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ _05438_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__nor2_1
X_11201_ _04264_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12181_ _05362_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nand2_1
X_11132_ _04211_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__xor2_4
X_11063_ _03589_ _03597_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__o21ai_4
X_10014_ net43 net39 net40 net42 VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11965_ _05124_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__or2_1
X_10916_ _03376_ _03378_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11896_ _05028_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__xor2_4
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10847_ _03896_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10778_ _03217_ _03219_ _03218_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12517_ _05130_ _05135_ _05481_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__a31o_4
X_12448_ _05651_ _05655_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12379_ _05562_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06940_ net96 VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06871_ _02394_ _06171_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__and3_1
X_08610_ _01508_ _01509_ _01496_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a21o_1
X_09590_ _01860_ _01867_ _01866_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__a21boi_1
X_08541_ _00874_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__xnor2_2
X_08472_ _01363_ _01372_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07423_ _00314_ _00325_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07354_ _00246_ _00255_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07285_ _06232_ _00187_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09024_ _01920_ _01921_ _01922_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09926_ _02266_ _02299_ _02298_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09857_ _02148_ _02149_ _02150_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__and3_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _02725_ _02738_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__xnor2_2
X_08808_ _01706_ _01707_ _01113_ net318 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__a211o_1
X_08739_ _01637_ _01638_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__nand3_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _04491_ _04526_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__a21o_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _03248_ _03312_ _03310_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a21o_2
X_11681_ _03881_ _04397_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__and2_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _03662_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__xor2_4
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10563_ _03577_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12302_ _05162_ _05157_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10494_ _03510_ _03511_ _03485_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12233_ _05410_ _05419_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12164_ _05342_ _05344_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__xor2_1
X_11115_ _04191_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__xor2_4
X_12095_ _05233_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xnor2_2
X_11046_ _03532_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11948_ _04974_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11879_ _05031_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07070_ net238 VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09711_ _02582_ _02583_ _02652_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__a211o_1
X_07972_ _03732_ net50 _00397_ _00872_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__and4_2
XFILLER_0_93_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06923_ _06197_ _06201_ _06235_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__and3_1
X_09642_ _02484_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__xnor2_4
X_06854_ _02536_ _04205_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__and2b_1
X_06785_ net237 VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__buf_4
X_09573_ _00200_ _00238_ _00703_ net88 VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08524_ _01379_ _00862_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08455_ _01353_ _01354_ _01174_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__a21o_1
X_08386_ _00747_ _00751_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__or2b_1
X_07406_ _00306_ _00307_ _00308_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07337_ net25 _06261_ _00239_ net24 VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07268_ net170 VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_4
X_09007_ net149 _01309_ _01904_ _01905_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__nand4_1
X_07199_ _04884_ _00102_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09909_ _02869_ _02870_ _02860_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__a21o_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ net272 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__inv_2
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _00872_ _01444_ _01434_ _02765_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _05878_ _05934_ _05948_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__o21ai_1
X_11733_ _04867_ _04871_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__xor2_4
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11664_ _00672_ _01835_ _04320_ _04321_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a31o_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10615_ _03013_ _03028_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__a21o_2
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11595_ net260 _04720_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__nor2_1
X_10546_ _02966_ _02975_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__a21o_2
XFILLER_0_121_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10477_ _02863_ _02865_ _02864_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12216_ _05401_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or2_4
XFILLER_0_102_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12147_ _01443_ _02799_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nand2_1
X_12078_ _05250_ _04866_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__or2_4
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11029_ _04098_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06570_ _02668_ _03612_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08240_ _00178_ _00625_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08171_ net1 _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07122_ _03425_ _05422_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07053_ _05958_ _06045_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07955_ _00854_ _00855_ _00398_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__a21o_1
X_06906_ _06219_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__nand2_1
X_09625_ _01874_ _01876_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nand2_1
X_07886_ _00740_ _00786_ _00787_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__and3_1
X_06837_ net124 VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__clkbuf_4
X_06768_ _05783_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__inv_2
X_09556_ _02454_ _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__xnor2_4
X_08507_ _05914_ _00822_ _01406_ _01407_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__a22o_1
X_06699_ _02822_ _03194_ _03183_ _05027_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a31o_2
X_09487_ _01763_ _01729_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__or2b_1
X_08438_ _01307_ _01337_ _01338_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__nor3_2
XFILLER_0_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08369_ _00679_ _00681_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11380_ _04474_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__xnor2_2
X_10400_ _02773_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__xor2_1
X_10331_ _03321_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10262_ _00291_ net153 _01288_ net142 VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__a22o_1
X_12001_ _05155_ _05156_ _05165_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a21o_1
X_10193_ _03179_ _03181_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12903_ clknet_1_1__leaf_clk _00027_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dfxtp_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _02174_ _06075_ _06076_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _05997_ _05928_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__a21oi_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _00343_ _03859_ _04404_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__and3_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12696_ _05915_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__nand2_1
Xinput13 data_in[110] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11647_ _04776_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput46 data_in[140] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput35 data_in[130] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 data_in[120] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11578_ _04701_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__xor2_4
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput68 data_in[160] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
Xinput79 data_in[170] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
Xinput57 data_in[150] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
X_10529_ _02931_ _02935_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07740_ net166 net161 net162 net165 VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07671_ _00571_ _00572_ _00528_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__o21a_1
X_06622_ _04117_ _04172_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__nand2_1
X_09410_ _02322_ _02323_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__nor2_1
X_09341_ _02236_ _02246_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06553_ _03359_ _03370_ _03403_ _03425_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09272_ net89 _01524_ _02170_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06484_ _02635_ _02646_ _02657_ _02668_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08223_ _01123_ _01124_ _00595_ _00597_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__o211a_1
X_08154_ _04862_ net36 net37 _03194_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08085_ net183 net182 _00058_ _00481_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__and4_1
X_07105_ _05411_ _06417_ _06418_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07036_ _02580_ _06347_ _06349_ _06346_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08987_ _01884_ _01885_ _01303_ _01305_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__o211a_1
X_07938_ _00838_ _00839_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__xnor2_1
X_07869_ _00298_ _00305_ _00304_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10880_ _00366_ _02694_ _02695_ _06383_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__a22o_1
X_09608_ _02538_ _02539_ _02516_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__o21a_1
X_09539_ _06130_ _01188_ _02464_ _04238_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ _05577_ _05579_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11501_ _04148_ _04149_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12481_ _05008_ _05691_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__a21oi_1
X_11432_ _04537_ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11363_ _04464_ _04465_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11294_ _01309_ _04389_ _04390_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__a21bo_1
X_10314_ _03126_ _03314_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__xor2_4
X_10245_ _02543_ _02571_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a21oi_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10176_ _03162_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12817_ _06018_ _06025_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ net265 _05983_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12679_ _05823_ _05824_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap302 _00569_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_1
XFILLER_0_25_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08910_ _06253_ _00200_ _01808_ _01809_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a22oi_1
X_09890_ _02814_ _02849_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__and3_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _01739_ _01740_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__xnor2_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _01670_ _01671_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__nand3_1
XFILLER_0_109_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07723_ _00623_ _00624_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__xnor2_2
X_07654_ _00553_ _00554_ _00555_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06605_ _03776_ _03985_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07585_ _00478_ _00487_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06536_ _02866_ _03238_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nand2_1
X_09324_ _01566_ _01574_ _01573_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__a21bo_1
X_06467_ net243 VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__buf_4
X_09255_ _01508_ _01510_ _02153_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08206_ _00971_ _00973_ _01105_ _01106_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09186_ _03732_ _01434_ _02083_ _02084_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__nand4_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08137_ _00513_ _01038_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08068_ _00967_ _00968_ _00909_ _00502_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_3_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07019_ _06331_ _06332_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__nand2_1
X_10030_ _04939_ net56 net67 _03095_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__a22o_1
Xinput236 data_in[81] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xinput203 data_in[51] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
Xinput214 data_in[61] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
Xinput225 data_in[71] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xinput247 data_in[91] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_2
X_11981_ _05130_ _05135_ _05128_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a21boi_2
X_10932_ _03991_ _03992_ _03406_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10863_ _03432_ _03516_ _03515_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__a21boi_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10794_ _03840_ _03841_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12602_ _05823_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12533_ _05493_ _05514_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _05666_ _05673_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12395_ _01410_ _01397_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_1
X_11415_ _03982_ _04012_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11346_ _03928_ _04445_ _04447_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_61_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11277_ _04370_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__xnor2_4
X_10228_ _03217_ _03218_ _03219_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__nand3_1
X_10159_ _06138_ net31 VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07370_ _02317_ _04238_ _06243_ _00270_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09040_ _01938_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09942_ _00047_ _00058_ _00489_ _00481_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09873_ net116 net108 net109 net115 VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__a22o_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _01722_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__xor2_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _01654_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__nor2_1
X_07706_ _00605_ _00606_ _00607_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__or3_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _01584_ _01585_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__a21bo_1
X_07637_ _00103_ _00539_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__nand2_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ _00468_ _00469_ _00034_ _00037_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09307_ _02202_ _02210_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06519_ _03053_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07499_ _05783_ _05805_ _06352_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09238_ _02135_ _02136_ _01486_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09169_ _02065_ _02066_ _02067_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__nand3_1
XFILLER_0_133_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11200_ _04265_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__xnor2_4
X_12180_ _04993_ _05361_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11131_ _03569_ _03657_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11062_ _03594_ _03596_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__or2b_1
X_10013_ _02984_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11964_ _04256_ _04717_ _05125_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__a21oi_1
X_10915_ _03960_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__xor2_2
X_11895_ _05041_ _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__xor2_4
XFILLER_0_129_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10846_ _03285_ _03898_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10777_ _03819_ _03821_ _03822_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12516_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12447_ _05651_ _05655_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12378_ _05577_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11329_ _04426_ _04428_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06870_ _04183_ _06184_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__xor2_1
X_08540_ _01439_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08471_ _01370_ _01371_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07422_ _00323_ _00324_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07353_ _00246_ _00255_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07284_ _00185_ _00186_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09023_ _01920_ _01921_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09925_ _02795_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__xnor2_4
X_09856_ _02796_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__xnor2_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _01113_ net318 _01706_ _01707_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__o211ai_4
X_09787_ _02730_ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__xnor2_2
X_06999_ _06178_ _04150_ _06312_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__a21o_1
X_08738_ _01055_ _01056_ _01057_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__a21bo_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08669_ _03337_ _01567_ _01568_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__nand4_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _03697_ _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__xnor2_2
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04812_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10631_ _02890_ _03044_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10562_ _03586_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12301_ _05166_ _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nand2_2
XFILLER_0_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12232_ _05410_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__or2_1
X_10493_ _03485_ _03510_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12163_ _04942_ _04963_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__a21o_1
X_11114_ _04192_ _04193_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__nor2_2
XFILLER_0_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12094_ _05265_ _05267_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__xor2_2
X_11045_ _00062_ _02215_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11947_ _05105_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11878_ _01002_ _01584_ _01562_ _02904_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10829_ _03287_ _03879_ _03880_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07971_ _03732_ _00397_ _00872_ net50 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__a22oi_1
X_09710_ _02650_ _02651_ _02584_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__o21a_1
X_06922_ _06197_ _06201_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09641_ _02575_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__xor2_4
X_06853_ _06133_ _06165_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__nand2_1
X_06784_ net246 VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__clkbuf_4
X_09572_ _02499_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__nor2_1
X_08523_ _01403_ _01423_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08454_ _01174_ _01353_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__nand3_1
X_07405_ _06175_ _06309_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__and2_1
X_08385_ _00808_ _00814_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07336_ net19 VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ net149 net146 _01904_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07267_ _06226_ _06234_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__nand2_1
X_07198_ _00099_ _00101_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09908_ _02860_ _02869_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__nand3_2
X_09839_ _02794_ _02190_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__or2_2
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12850_ _06091_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__clkbuf_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _01444_ _01434_ _02765_ _00872_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a22oi_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12781_ _05543_ _05774_ _05937_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__and3_2
X_11732_ _04869_ _04870_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__nor2_2
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _00703_ _01251_ _01835_ _01858_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__nand4_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10614_ _03026_ _03027_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11594_ net260 _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__and2_1
X_10545_ _02974_ _02973_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10476_ _03489_ _03490_ _03492_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nand3_1
X_12215_ _05395_ _05399_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12146_ _04553_ _04980_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__nand2_1
X_12077_ net216 VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__inv_2
X_11028_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08170_ net45 VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07121_ _06414_ _06432_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07052_ _06364_ _06365_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07954_ _00398_ _00854_ _00855_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07885_ _00784_ _00785_ _00741_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__a21o_1
X_06905_ net269 _04666_ _04688_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a21boi_1
X_06836_ net132 VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__buf_2
X_09624_ _02548_ _02557_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__xnor2_2
X_06767_ _03732_ _03743_ _02580_ _05761_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__and4_1
X_09555_ _02455_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xnor2_4
X_08506_ _05882_ _06375_ _06368_ net2 VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__nand4_2
X_06698_ _02844_ _03172_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__and2_1
X_09486_ _00166_ _02407_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08437_ _01335_ _01336_ _01308_ _00780_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08368_ _01267_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07319_ _00198_ _00199_ _00220_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__nor3_1
XFILLER_0_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08299_ _01178_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__xnor2_2
X_10330_ _03323_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10261_ net142 net143 net154 VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12000_ _05163_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__xor2_1
X_10192_ _06159_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ clknet_1_1__leaf_clk _00026_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ _06071_ _06074_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__nand2_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12764_ _05998_ _06000_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__xnor2_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _04394_ _04396_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12695_ _05916_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11646_ _00647_ _02498_ _04775_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__and3_1
Xinput36 data_in[131] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
Xinput25 data_in[121] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput14 data_in[111] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_0_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11577_ _04092_ _04214_ _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput69 data_in[161] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput58 data_in[151] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xinput47 data_in[141] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
X_10528_ _03530_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__xor2_4
XFILLER_0_122_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10459_ _03473_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
X_12129_ _04949_ _04951_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__and2b_1
X_07670_ _00528_ _00571_ _00572_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__nor3_1
X_06621_ _04117_ _04172_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09340_ _02244_ _02245_ _02237_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06552_ _03414_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__inv_2
X_09271_ net100 net111 _00453_ _00953_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand4_2
X_06483_ net68 VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__buf_2
X_08222_ _01121_ _01122_ _00612_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08153_ _04906_ _00097_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08084_ _02734_ _00985_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__nand2_1
X_07104_ net104 net103 _05444_ _06416_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__nand4_1
XFILLER_0_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07035_ _06345_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08986_ _01303_ _01305_ _01884_ _01885_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__a211oi_4
X_07937_ _00371_ _00372_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__nand2_1
X_07868_ _00767_ _00768_ _00760_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06819_ net96 VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__clkbuf_4
X_09607_ _02516_ _02538_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__nor3_1
X_07799_ _00699_ _00698_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09538_ net164 VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ _04099_ _04617_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09469_ _01764_ _02387_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nand3_2
X_12480_ _01563_ _01524_ _02215_ _03499_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11431_ _04540_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11362_ _03948_ _03950_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10313_ _03129_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11293_ net153 net146 _01288_ _00774_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a22o_1
X_10244_ _02544_ _02570_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__and2_1
X_10175_ net26 net27 net21 net22 VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nand4_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12816_ _06031_ _06033_ _06029_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12747_ net265 _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__nand2_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _05821_ _05831_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11629_ _04735_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08840_ _06127_ _00617_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__nand2_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _01078_ _01080_ _01079_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__a21bo_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ _00172_ _00175_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__nand2_1
X_07653_ _00553_ _00554_ _00555_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__nand3_2
X_06604_ _03776_ _03985_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09323_ _02225_ _02226_ _02217_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a21o_1
X_07584_ _00061_ _00486_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__xnor2_1
X_06535_ _03227_ net226 net227 VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06466_ net252 VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09254_ _02151_ _02152_ _02140_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09185_ _03732_ _01434_ _02083_ _02084_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__a22o_1
X_08205_ _00971_ _00973_ _01105_ _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__nor4_2
XFILLER_0_28_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08136_ net226 _03260_ _00507_ _01034_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08067_ _00909_ _00502_ _00967_ _00968_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_31_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07018_ _06302_ _06303_ _06330_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__or3_2
XFILLER_0_3_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput204 data_in[52] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
Xinput215 data_in[62] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
Xinput226 data_in[72] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_2
Xinput248 data_in[92] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
Xinput237 data_in[82] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_4
X_08969_ _01866_ _01867_ _01860_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__a21oi_1
X_11980_ _05143_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10931_ _03406_ _03991_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10862_ _03422_ _03424_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10793_ _03837_ _03839_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__nand2_1
X_12601_ _05649_ _05659_ _05647_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ _05515_ _05491_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12463_ _05671_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11414_ _04011_ _03983_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12394_ _05299_ _05300_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11345_ _04445_ _04447_ _03928_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11276_ _03814_ _03836_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a21o_2
X_10227_ _03217_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__a21o_1
X_10158_ _03142_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nand2_1
X_10089_ _03067_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09941_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09872_ net114 net109 _02166_ _02165_ net110 VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__a32o_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _01129_ _01130_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _02800_ net41 _01652_ _01653_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _00605_ _00606_ _00607_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__o21ai_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08685_ net192 net187 net188 net191 VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07636_ _00531_ _00538_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__xnor2_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07567_ _00034_ _00037_ _00468_ _00469_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a211oi_2
X_09306_ _02208_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__or2b_1
X_06518_ _02185_ _03031_ _03042_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07498_ _00396_ _00400_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__xnor2_1
X_09237_ _01486_ _02135_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06449_ _02196_ _02207_ _02262_ _02284_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__nand4_2
X_09168_ _02065_ _02066_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09099_ _01370_ _01996_ _01997_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08119_ _00515_ _00524_ _00514_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11130_ _03653_ _03655_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11061_ _04094_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__xnor2_4
X_10012_ _04906_ net48 VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11963_ _04714_ _04716_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10914_ _03971_ _03973_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__xnor2_2
X_11894_ _05047_ _05048_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__nand2_2
X_10845_ _03297_ _03298_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10776_ _03819_ _03821_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12515_ _05128_ _05478_ _05480_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12446_ _05653_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__xnor2_1
X_12377_ _05236_ _05264_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11328_ _04426_ _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11259_ _00210_ _00677_ net137 net138 VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__and4_1
X_08470_ _01364_ _01369_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__nor2_1
X_07421_ _06315_ _00322_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07352_ _06265_ _00254_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07283_ _00184_ _00183_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__and2b_1
X_09022_ net211 net204 VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09924_ _02886_ _02887_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__or2b_2
X_09855_ _02810_ _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__or2b_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _01355_ _01356_ _01704_ _01705_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__a22o_1
X_09786_ _02735_ _02736_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__xnor2_2
X_06998_ _02383_ _04139_ _06177_ _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__nand4_2
X_08737_ net36 _00097_ _01635_ _01636_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08668_ net184 _00047_ _00058_ _00480_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__nand4_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _00088_ _00521_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _03041_ _03043_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__nor2_1
X_08599_ _05444_ net106 net116 net107 VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ _03583_ _03584_ _03585_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10492_ _03508_ _03509_ _02878_ _03486_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _05154_ _05168_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12231_ _05414_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12162_ _04940_ _04964_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__and2_1
X_11113_ _00549_ _00550_ net56 _03006_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__and4_2
X_12093_ _04844_ _04879_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__a21oi_2
X_11044_ _05202_ _01563_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11946_ _04599_ _04700_ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__o21a_2
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11877_ _01584_ _01562_ _02904_ _01002_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a22oi_1
X_10828_ _06362_ _03859_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10759_ _03796_ _03802_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12429_ _05620_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07970_ net64 VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06921_ _06226_ _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__xnor2_1
X_09640_ _01890_ _01892_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__nand2_2
X_06852_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__inv_2
X_06783_ _05893_ _05947_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09571_ _04292_ _04446_ net102 _02498_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__and4_2
X_08522_ _01421_ _01422_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08453_ _01351_ _01352_ _00903_ _00905_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__a211o_1
X_07404_ _00304_ _00305_ _00298_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08384_ _00782_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07335_ net98 VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07266_ _00152_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09005_ net199 net216 net147 net148 VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07197_ _02822_ _00097_ _00098_ _00100_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09907_ _02867_ _02868_ _02861_ _02862_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__a211o_1
X_09838_ _02188_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__inv_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _02714_ _02715_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nand3_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04945_ _04542_ _04546_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__a21o_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12780_ _05757_ _05962_ _05960_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__a21oi_4
X_11731_ _00810_ _03859_ _04408_ _04868_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11662_ _01251_ _01835_ _01858_ _00703_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__a22o_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10613_ _03629_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__xor2_4
XFILLER_0_107_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11593_ _04251_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10544_ _03521_ _03567_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10475_ _03489_ _03490_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__a21o_1
X_12214_ _05395_ _05399_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__nor2_1
X_12145_ _03999_ _04511_ _04958_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__a31o_2
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12076_ _02626_ _01986_ _03859_ _01365_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a22oi_1
X_11027_ _00047_ net186 net197 net198 VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__and4_2
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11929_ _05086_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07120_ _06433_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07051_ _02503_ _03886_ _06034_ _02448_ _06362_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07953_ _00848_ _00849_ _00851_ _00853_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__a22o_1
X_07884_ _00741_ _00784_ _00785_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__nand3_2
X_06904_ net278 _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__xnor2_1
X_09623_ _02555_ _02556_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__and2b_1
X_06835_ _06148_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06766_ _03732_ _03743_ _02580_ _05761_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a22o_1
X_09554_ _02457_ _02480_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__xnor2_4
X_06697_ _04895_ _05005_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__xnor2_4
X_08505_ net255 net9 net2 net8 VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ _02404_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__xor2_1
X_08436_ _01308_ _00780_ _01335_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08367_ _06151_ _00210_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07318_ _00198_ _00199_ _00220_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08298_ _00651_ _01198_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__xor2_2
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07249_ _00149_ _00150_ _00151_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10260_ _02612_ _02619_ _02618_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10191_ net102 VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__clkbuf_4
X_12901_ clknet_1_1__leaf_clk _00025_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dfxtp_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12832_ _06071_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__or2_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12763_ _05999_ _05920_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__xnor2_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _03868_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _05923_ _05924_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11645_ _00647_ _02498_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput37 data_in[132] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
Xinput26 data_in[122] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_4
Xinput15 data_in[112] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11576_ _04211_ _04213_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 data_in[152] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
Xinput48 data_in[142] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10527_ _03548_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10458_ _03471_ _03472_ _02823_ _02825_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10389_ _06343_ net65 _03396_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__a22o_1
X_12128_ _00879_ _03967_ _04923_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__and3_1
X_12059_ _04831_ _04833_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__and2b_1
X_06620_ _02394_ _04150_ _04161_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06551_ _03381_ net167 _03392_ _02745_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06482_ net76 VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__clkbuf_4
X_09270_ net111 net177 net178 net100 VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__a22o_1
X_08221_ _00612_ _01121_ _01122_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__nor3_1
XFILLER_0_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08152_ _01052_ _01053_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08083_ net134 VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_4
X_07103_ net104 _05444_ _06416_ net103 VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__a22o_1
X_07034_ _06345_ _06346_ net50 _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__and4b_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _01882_ _01883_ _01870_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__a21oi_2
X_07936_ _00836_ _00837_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__or2_1
X_07867_ _00760_ _00767_ _00768_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09606_ _02535_ _02537_ _02517_ _02518_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__a211oi_1
X_07798_ _00698_ _00699_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06818_ _04490_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09537_ _01220_ _01824_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__a21bo_2
X_06749_ _03623_ _05575_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09468_ _02385_ _02386_ _01765_ _01766_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__a211o_1
X_09399_ net43 net38 net39 net42 VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__a22o_1
X_08419_ _02459_ net215 VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11430_ _01487_ _00937_ _04030_ _04028_ _02799_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11361_ _04462_ _04463_ _03965_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10312_ _03248_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11292_ _00774_ net153 _01288_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10243_ _03207_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10174_ net27 net21 net22 net26 VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12815_ _06005_ _06013_ _06003_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12746_ _05977_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12677_ _05905_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11628_ _04736_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11559_ _04675_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap304 _02233_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _01668_ _01669_ _01665_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__a21o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07721_ _00620_ _00622_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__nand2_1
X_07652_ _00111_ _00113_ _00112_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__a21bo_1
X_07583_ _00484_ _00485_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__and2b_1
X_06603_ _03963_ _03974_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__nor2_1
X_06534_ net218 VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__buf_2
XFILLER_0_87_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09322_ _02217_ _02225_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06465_ net6 VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__clkbuf_4
X_09253_ _02140_ _02151_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__and3_2
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09184_ _05750_ net53 _00397_ _00872_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__nand4_2
XFILLER_0_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08204_ net294 _01104_ _00575_ _00577_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08135_ _00508_ _01036_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08066_ _00949_ _00950_ _00966_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07017_ _06302_ _06303_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput216 data_in[63] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_4
Xinput205 data_in[53] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_4
Xinput227 data_in[73] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_2
Xinput249 data_in[93] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_2
Xinput238 data_in[83] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_4
X_08968_ _01860_ _01866_ _01867_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__and3_1
X_07919_ net11 VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_4
X_08899_ _01772_ _01243_ _01797_ _01798_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__o211ai_4
X_10930_ _00387_ net65 _03989_ _03990_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10861_ _03385_ _03426_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__or2b_1
X_12600_ _05821_ _05822_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__and2_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _03837_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12531_ _05730_ _05733_ _05727_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__a21oi_4
X_12462_ _05420_ _05424_ _05670_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11413_ _04493_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__xnor2_2
X_12393_ _05594_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11344_ _03938_ _03942_ _04444_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__or3_1
X_11275_ _03815_ _03835_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10226_ net126 net136 VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__and2_1
X_10157_ net18 net19 _00647_ _01181_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10088_ net284 _03066_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12729_ _05957_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09940_ net183 net184 net197 net198 VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__and4_2
X_09871_ _02143_ _02145_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ net281 _01128_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _02800_ _01652_ _01653_ net41 VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__a22oi_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ _00163_ _00164_ _00162_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08684_ net191 net192 _01002_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07635_ _00536_ _00537_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__xor2_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ _00466_ _00467_ _00075_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09305_ _02205_ _02206_ _01565_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06517_ net258 _03009_ _03020_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07497_ _00398_ _00399_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09236_ net103 _02132_ _02133_ _02134_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__nand4_1
XFILLER_0_106_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06448_ _02273_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__inv_2
X_09167_ net59 net58 VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09098_ _01996_ _01997_ _01370_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__a21o_1
X_08118_ _00974_ _00975_ _01018_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08049_ _00061_ _00486_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11060_ _04097_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__xnor2_4
X_10011_ _02982_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11962_ _04729_ _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__xor2_1
X_10913_ _03364_ _03375_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a21oi_2
X_11893_ _04623_ _05046_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10844_ _03297_ _03298_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10775_ net127 net136 VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__and2_1
X_12514_ _05727_ _05728_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__nor2_2
X_12445_ _05068_ _04154_ _02329_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__and3b_1
X_12376_ _05238_ _05263_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11327_ _03850_ _03905_ _04427_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_105_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11258_ _00677_ net137 net138 _00210_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10209_ _03188_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__xnor2_1
X_11189_ _03717_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__xnor2_1
X_07420_ _06315_ _00322_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07351_ _00252_ _00253_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07282_ _00183_ _00184_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09021_ _04106_ _06173_ net205 net206 VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__nand4_2
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09923_ _02884_ _02885_ _02259_ _02261_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09854_ _02808_ _02809_ _02797_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__a21o_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _01355_ _01356_ _01704_ _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nand4_2
X_09785_ _02042_ _02044_ _02041_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__o21bai_2
X_06997_ net142 VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__clkbuf_4
X_08736_ _00107_ _00097_ _01635_ _01636_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__nand4_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _00047_ _00989_ _00480_ net184 VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__a22o_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _00517_ _00520_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08598_ net106 net116 net107 net115 VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07549_ _00430_ _00451_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__xor2_2
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10560_ _03583_ _03584_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09219_ _01490_ _01492_ _02117_ _02118_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a211o_1
X_10491_ _02878_ _03486_ _03508_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12230_ _05415_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__xor2_2
X_12161_ _05320_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__xnor2_2
X_11112_ _00550_ _01652_ _03006_ _00549_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__a22oi_1
X_12092_ _04846_ _04878_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nor2_1
X_11043_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11945_ _04696_ _04698_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11876_ _04609_ _04613_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__nand2_1
X_10827_ _06362_ _02626_ _03288_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__and3_1
X_10758_ _03796_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10689_ _03104_ _03110_ _03725_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nor3_1
X_12428_ _05621_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12359_ _05226_ _05540_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06920_ _06232_ _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nor2_1
X_06851_ _06133_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__nor2_1
X_06782_ _05904_ _05925_ _05936_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__or3_2
XFILLER_0_89_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09570_ _04292_ net102 _02498_ _04446_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__a22oi_2
X_08521_ _01418_ _01419_ _01420_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08452_ _00903_ _00905_ _01351_ _01352_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__o211ai_2
X_07403_ _00298_ _00304_ _00305_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08383_ _01283_ _00788_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07334_ _00235_ _00236_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07265_ _06211_ _00156_ _00157_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09004_ net199 net148 net216 net147 VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__nand4_2
XFILLER_0_131_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07196_ _00096_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2 _01111_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09906_ _02861_ _02862_ _02867_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o211ai_2
X_09837_ _02667_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__xor2_4
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _02029_ _02027_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__o21a_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _01053_ _01618_ _01619_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__and3_1
X_09699_ _02638_ _02639_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__and3_1
X_11730_ _04408_ _04868_ _00810_ _03859_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__o211a_2
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _00200_ _03180_ _04328_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__nand3_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10612_ _03640_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11592_ _04253_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10543_ _03523_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10474_ net111 net180 VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12213_ _05396_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__xor2_1
X_12144_ _04952_ _04959_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12075_ _04867_ _04869_ _04870_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__or3_1
X_11026_ _00489_ net197 net198 _00049_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11928_ _01068_ _04154_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11859_ _05009_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07050_ _03897_ _06012_ _06023_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__or4_2
XFILLER_0_82_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07952_ _00848_ _00849_ _00851_ _00853_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__nand4_2
X_07883_ _00782_ _00783_ _00755_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__o21ai_2
X_06903_ _06216_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__xor2_2
XFILLER_0_128_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09622_ _02553_ _02554_ _02549_ _02550_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__a211o_1
X_06834_ _06137_ _06147_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09553_ _02458_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__xnor2_4
X_08504_ _00355_ _01404_ _00854_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a21bo_1
X_06765_ net61 VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06696_ _03150_ _04994_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__xor2_4
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _01721_ _01724_ _01720_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__a21o_1
X_08435_ _01333_ _01334_ _01316_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__o21a_1
X_08366_ _01264_ _01265_ _01266_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07317_ _06323_ _00219_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08297_ _01179_ _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07248_ _00149_ _00150_ _00151_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__or3_2
XFILLER_0_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07179_ _03260_ _04752_ _00082_ _00080_ _02855_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10190_ _03177_ _03178_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__xnor2_1
X_12900_ clknet_1_1__leaf_clk _00024_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dfxtp_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12831_ _05987_ _05993_ _06047_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__a31o_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12762_ _05905_ _05906_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or2_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _04440_ _04454_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a21o_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12693_ _05917_ _05918_ _05922_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _01217_ _01181_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 data_in[123] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_4
Xinput16 data_in[113] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11575_ _04599_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput49 data_in[143] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
Xinput38 data_in[133] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
X_10526_ _03544_ _03545_ _03547_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10457_ _02823_ _02825_ _03471_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10388_ net54 net63 net55 net64 VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand4_2
X_12127_ _05303_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__nor2_1
X_12058_ _05212_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__xor2_4
X_11009_ _04076_ _04077_ _04061_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06550_ _03381_ _02734_ _03392_ _02745_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06481_ net103 VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08220_ _01119_ _01120_ _00591_ _00593_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08151_ _03084_ net32 _00530_ _01051_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08082_ _00982_ _00983_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__or2_1
X_07102_ net116 VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__clkbuf_4
X_07033_ net62 VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08984_ _01870_ _01882_ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07935_ _05969_ _06384_ _00833_ _00835_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__and4_2
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07866_ _00765_ _00766_ _00761_ _00762_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__a211o_1
X_09605_ _02517_ _02518_ _02535_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__o211a_1
X_07797_ _00248_ _00251_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__nand2_1
X_06817_ _06129_ _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__xor2_2
X_09536_ _01825_ _01819_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__or2b_1
X_06748_ _05477_ _05564_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09467_ _01765_ _01766_ _02385_ _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__o211ai_2
X_08418_ _01317_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__nor2_1
X_06679_ _02866_ _04741_ _04807_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09398_ _00107_ _00097_ _01635_ _01636_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08349_ net137 VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11360_ _03965_ _04462_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_6_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10311_ _03310_ _03311_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11291_ _03921_ _03935_ _04387_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__a21o_2
XFILLER_0_30_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10242_ _03209_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10173_ _02542_ _02574_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12814_ _06052_ _06054_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__xnor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _05730_ _05733_ _05899_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _05436_ _05692_ _05828_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11627_ _04737_ _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__xor2_4
X_11558_ _04680_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap305 _02091_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_1
X_10509_ _03525_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__xor2_4
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11489_ _00481_ _01567_ net188 _02239_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _00621_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__inv_2
X_07651_ _00551_ _00552_ _00548_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__a21o_1
X_07582_ _02734_ _00479_ _00482_ _00483_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a22o_1
X_06602_ _03930_ _03952_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__and2_1
X_06533_ _03183_ _03205_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__xnor2_4
X_09321_ _02223_ _02224_ _02219_ _02220_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06464_ net199 VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_4
X_09252_ _02148_ _02149_ _02150_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09183_ net53 net63 net64 net52 VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08203_ _00575_ _00577_ net294 _01104_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_50_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08134_ _02855_ _03260_ _00507_ _01034_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__nand4_1
XFILLER_0_16_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08065_ _00949_ _00950_ _00966_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07016_ _06328_ _06329_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput217 data_in[64] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_2
Xinput206 data_in[54] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_4
Xinput228 data_in[74] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_4
Xinput239 data_in[84] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
X_08967_ _01863_ _01864_ _01865_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__a21o_1
X_07918_ _00365_ _00378_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__or2_1
X_08898_ _01795_ _01796_ _01773_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__a21bo_1
X_07849_ _00747_ _00748_ net139 _00749_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__or4bb_1
X_10860_ _03740_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xor2_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09519_ _02440_ _02441_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10791_ _03207_ _03236_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__a21oi_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12530_ _05746_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12461_ _05420_ _05424_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11412_ _04495_ _04520_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12392_ _05285_ _05593_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11343_ _03938_ _03942_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__o21ai_2
X_11274_ _04349_ _04368_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10225_ _06283_ _00201_ _00677_ net128 VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nand4_1
X_10156_ net19 net29 net30 net18 VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10087_ net284 _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10989_ _04055_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12728_ _05757_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__xor2_4
X_12659_ _05710_ _05712_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09870_ _02818_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__xnor2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _01720_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ net39 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_4
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ net188 VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_4
X_07703_ _00601_ _00604_ net280 VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__a21oi_1
X_07634_ _00096_ _00099_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07565_ _00075_ _00466_ _00467_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__and3_1
X_07496_ _02580_ _00397_ _06345_ _06348_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__a211oi_1
X_09304_ _01565_ _02205_ _02206_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06516_ _03009_ _03020_ net258 VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06447_ _02218_ _02229_ _02240_ _02251_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__and4_2
X_09235_ net103 _02132_ _02133_ _02134_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09166_ net69 net68 _01443_ _02064_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__nand4_1
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09097_ _01994_ _01995_ _01985_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08117_ _00974_ _00975_ _01018_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08048_ _00935_ _00936_ _00948_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ net36 net37 net46 net47 VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__and4_1
X_09999_ _02969_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__or2b_1
X_11961_ _05120_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__xnor2_1
X_10912_ _03365_ _03374_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__and2_1
X_11892_ _04623_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10843_ _03883_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__xor2_2
X_10774_ net133 net135 net128 net129 VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__nand4_1
XFILLER_0_109_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12513_ _05486_ _05488_ _05726_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12444_ _03580_ _04123_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12375_ _05563_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11326_ _03852_ _03904_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11257_ _06311_ _02592_ _03862_ _03861_ _00749_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10208_ _03197_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__and2b_1
X_11188_ _04273_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__nor2_1
X_10139_ _03086_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07350_ _00249_ _00251_ _06263_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09020_ _06172_ net205 net206 net209 VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07281_ _06252_ _06298_ _06297_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09922_ _02259_ _02261_ _02884_ _02885_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09853_ _02797_ _02808_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__and3_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _02732_ _02733_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__nor2_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _01702_ _01703_ _01109_ net290 VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__a211o_1
X_08735_ _03194_ _04862_ _00543_ _01068_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__nand4_2
X_06996_ _06175_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__xnor2_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08666_ net196 VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07617_ _04741_ _00518_ _00519_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__a21bo_1
X_08597_ net113 net114 _00454_ _00956_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07548_ _00449_ _00450_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__xor2_2
XFILLER_0_49_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07479_ _00379_ _00380_ _00349_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09218_ _05498_ _00937_ _02115_ _02116_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__and4_1
X_10490_ _03506_ _03507_ _02873_ _02875_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09149_ _02034_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12160_ _05339_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__nor2_1
X_11111_ _03630_ _03632_ _03631_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a21bo_2
X_12091_ _05236_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11042_ _04111_ _04112_ _04113_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11944_ _05024_ _05103_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11875_ _04607_ _04608_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__nand2_1
X_10826_ _03876_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10757_ _03797_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10688_ _03104_ _03110_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12427_ _05632_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12358_ _05546_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__xnor2_1
X_11309_ _00297_ net214 net206 net207 VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12289_ net262 _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06850_ _04523_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06781_ _05914_ _03787_ net252 VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__and3b_1
XFILLER_0_117_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08520_ _01418_ _01419_ _01420_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__and3_1
X_08451_ _01349_ _01350_ _01282_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07402_ _00301_ _00302_ _00303_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08382_ _00786_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07333_ _00226_ _00234_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ _00165_ _00167_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ _01317_ _01320_ _01318_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07195_ _00096_ _00097_ net32 _00098_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__and4b_1
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09905_ _02863_ _02864_ _02865_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09836_ _02669_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__xnor2_4
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _02022_ _02023_ _02024_ _02025_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a211o_1
X_06979_ _06272_ _06291_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__or2_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _01917_ _01926_ _01925_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__a21bo_1
X_08718_ net226 net227 _01034_ _01617_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__nand4_2
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _01547_ _01548_ _01467_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__o21a_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _04327_ _04326_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__or2b_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _03018_ _03025_ _03641_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__a21oi_2
X_11591_ _04256_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10542_ _03551_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12212_ _04664_ _05059_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a21bo_1
X_10473_ _00479_ net177 net134 net178 VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12143_ _04985_ _05000_ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__o21a_1
X_12074_ _04869_ _05245_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__xnor2_2
X_11025_ _03571_ _03599_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a21o_2
XFILLER_0_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11927_ _04679_ _04681_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__nor2_1
X_11858_ _04572_ _04573_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10809_ net216 VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__clkbuf_4
X_11789_ _04481_ _04484_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07951_ _00355_ _00852_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06902_ _03073_ _04622_ _04633_ _04655_ _02350_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07882_ _00755_ _00782_ _00783_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__or3_4
X_09621_ _02549_ _02550_ _02553_ _02554_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__o211a_1
X_06833_ _06137_ _06147_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__nand2_1
X_06764_ net52 VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__clkbuf_4
X_09552_ _02461_ _02478_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__xor2_4
X_08503_ _00852_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__inv_2
X_06695_ _04917_ _04983_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__xnor2_4
X_09483_ _02402_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__or2b_1
X_08434_ _01316_ _01333_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__nor3_2
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08365_ net131 net127 net128 net130 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07316_ _00207_ _00218_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _00648_ _01196_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__xor2_2
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07247_ _06125_ _06203_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07178_ _03227_ _02855_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09819_ net69 _05498_ net83 net84 VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__and4_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _06072_ _06044_ _06046_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__o21ba_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12761_ _05821_ _05831_ _05907_ _05909_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__o22a_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04441_ _04453_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__nor2_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _05917_ _05918_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11643_ _04332_ _04334_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__a21oi_2
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 data_in[124] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput17 data_in[114] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
X_11574_ _04696_ _04698_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 data_in[134] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_0_134_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10525_ _03544_ _03545_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__and3_1
X_10456_ _03467_ _03468_ _03470_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10387_ net63 net55 net64 net54 VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__a22o_1
X_12126_ _05296_ _05302_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__and2_1
X_12057_ _05226_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11008_ _04061_ _04076_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06480_ net113 VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08150_ _03084_ _00530_ _01051_ _02822_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_74_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07101_ _05477_ _05531_ _05553_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08081_ _00981_ _00976_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07032_ net60 net52 net61 net51 VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08983_ _01880_ _01881_ _01871_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__a21o_1
X_07934_ _05969_ _06384_ _00833_ _00835_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07865_ _00761_ _00762_ _00765_ _00766_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__o211ai_2
X_09604_ _02533_ _02534_ _02520_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07796_ _00241_ _00697_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__xnor2_1
X_06816_ _02328_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06747_ _05531_ _05553_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__nor2_1
X_09535_ _01781_ _01782_ _01791_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o31ai_4
X_06678_ _04763_ _04796_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09466_ _02382_ _02384_ _01973_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__a21o_1
X_08417_ net200 _06077_ net213 net214 VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09397_ _03194_ _04862_ _00543_ _01068_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08348_ _00320_ _00753_ _00752_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08279_ _00241_ _00697_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11290_ _03922_ _03934_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__and2_1
X_10310_ _03308_ _03309_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ _03225_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__xnor2_2
X_10172_ _01886_ _01888_ _02572_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__o21ai_1
X_12813_ _06020_ _06022_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _05727_ _05978_ _05979_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05357_ _05844_ _05842_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11626_ _04753_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__nand2_2
XFILLER_0_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11557_ _04679_ _01629_ _01068_ _04676_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__and4b_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap306 _01091_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__buf_1
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10508_ _02906_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__xor2_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11488_ _01567_ _01584_ _02239_ _00481_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10439_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _05278_ _05280_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__a21o_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07650_ _00548_ _00551_ _00552_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__nand3_1
X_07581_ _02734_ _00479_ _00482_ _00483_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__and4_1
X_06601_ _03930_ _03952_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nor2_1
X_06532_ _02822_ _03194_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09320_ _02219_ _02220_ _02223_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09251_ _02148_ _02149_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06463_ net208 VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08202_ _01019_ _01020_ _01101_ _01102_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__o22a_2
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09182_ _06343_ _06347_ _01450_ _01449_ _00879_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08133_ _03260_ _00507_ _01034_ _02855_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08064_ _00461_ _00965_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__xnor2_1
X_07015_ _04183_ _06184_ _06186_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_113_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput218 data_in[65] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_2
Xinput207 data_in[55] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_2
Xinput229 data_in[75] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_4
X_08966_ _01863_ _01864_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__nand3_1
X_07917_ _06380_ _00364_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__nand2_1
X_08897_ _01773_ _01795_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__nand3b_2
X_07848_ _00747_ _00748_ _02394_ _00749_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07779_ _00678_ _00679_ net132 _06274_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__and4bb_1
X_09518_ _02440_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__nor2_1
X_10790_ _03209_ _03235_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__and2b_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _02302_ _02365_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__and3_2
XFILLER_0_94_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12460_ _05668_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12391_ _05285_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ _04497_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11342_ _04442_ _04443_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11273_ _04350_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10224_ net135 net127 net128 net133 VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10155_ _06130_ _02464_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10086_ _03061_ _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10988_ _03476_ _03465_ _03464_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12727_ _05960_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__and2b_2
X_12658_ _05815_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11609_ _04374_ _04375_ _04377_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_53_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12589_ _05807_ _05809_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ net282 _01719_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ net56 VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__buf_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ _02866_ _01023_ _01031_ _01030_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__a31o_1
X_07702_ net280 _00601_ _00604_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__and3_1
X_07633_ _00532_ _00535_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07564_ _00452_ _00465_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07495_ _06345_ _06348_ _02580_ _00397_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__o211a_1
X_09303_ net176 _00479_ _02203_ _02204_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06515_ _02987_ _02998_ _02437_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06446_ _02218_ _02229_ _02240_ _02251_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09234_ net104 net105 net118 net119 VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__nand4_2
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09165_ net69 net83 _02064_ net68 VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08116_ _00526_ _01017_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09096_ _01985_ _01994_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08047_ _00935_ _00936_ _00948_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_09998_ _03084_ net49 net225 net227 VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__a22o_1
X_08949_ _01817_ _01818_ _01848_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nor3b_1
X_11960_ _04293_ _04713_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__a21oi_1
X_10911_ _03961_ _03970_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__xnor2_2
X_11891_ _05043_ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10842_ _03892_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10773_ net135 net128 net129 net133 VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12512_ _05486_ _05488_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12443_ _01629_ _02329_ _05398_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12374_ _05565_ _05574_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11325_ _04382_ _04425_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__xnor2_1
X_11256_ _03858_ _03874_ _03873_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _02555_ _03189_ _03196_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__or3_1
X_11187_ _04269_ _04271_ _04272_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a21oi_1
X_10138_ _03089_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__xnor2_4
X_10069_ _02793_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07280_ net303 _00182_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09921_ _02851_ _02852_ _02882_ _02883_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09852_ _02806_ _02807_ _02798_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__a21o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ net51 _03798_ net66 net5 VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__and4_2
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _01109_ net290 _01702_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__o211ai_4
X_08734_ net43 net37 net38 net42 VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__a22o_1
X_06995_ _06305_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _01564_ _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nor2_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07616_ net219 net228 net229 net218 VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__a22o_1
X_08596_ _00922_ _00924_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__nand2_1
X_07547_ _06421_ _06429_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07478_ _00349_ _00379_ _00380_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__or3_2
XFILLER_0_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _05498_ _00937_ _02115_ _02116_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09148_ _02035_ _02047_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__xor2_2
XFILLER_0_91_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09079_ _01467_ _01547_ _01548_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _04188_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__or2b_2
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12090_ _05238_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__xor2_2
X_11041_ _04111_ _04112_ _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11943_ _05100_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__xor2_2
X_11874_ _04636_ _04656_ _04653_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a21o_2
XFILLER_0_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10825_ _03873_ _03874_ _03858_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10756_ _03212_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10687_ _03723_ _03724_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12426_ _05362_ _05365_ _05631_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12357_ _05555_ _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11308_ _00757_ _01365_ _01986_ _00297_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12288_ _05144_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__xnor2_2
X_11239_ _06284_ _03180_ _03788_ _03785_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a31o_1
X_06780_ _03820_ _03798_ _05914_ _02470_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08450_ _01282_ _01349_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07401_ _00301_ _00302_ _00303_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__and3_1
X_08381_ _01201_ _01281_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07332_ _00226_ _00234_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07263_ _00162_ _00163_ _00164_ _00166_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__a31o_1
X_07194_ net42 net35 net43 net33 VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__a22o_1
X_09002_ _00842_ _01374_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09904_ _02863_ _02864_ _02865_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__a21o_1
X_09835_ _02749_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__xnor2_4
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _02711_ _02713_ _02705_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a21o_1
X_06978_ _06272_ _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__nand2_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _02636_ _02637_ _02628_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__a21o_1
X_08717_ net227 _01034_ _01617_ net226 VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a22o_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _01467_ _01547_ _01548_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__nor3_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _00943_ _00941_ _00942_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ _03023_ _03024_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11590_ _04714_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10541_ _03562_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12211_ _04659_ _05058_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10472_ net177 net134 net178 net123 VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12142_ _04996_ _04999_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__or2b_1
X_12073_ _05243_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11024_ _03572_ _03598_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11926_ _00543_ _04154_ _04648_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11857_ _05007_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10808_ _03269_ _03272_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11788_ _04922_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10739_ _03780_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12409_ _05305_ _05311_ _05310_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07950_ net6 net7 net2 net3 VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__and4_2
XFILLER_0_121_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06901_ _06214_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__and2_1
X_07881_ _00780_ _00781_ _00756_ _00311_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09620_ _06274_ _00665_ _02551_ _02552_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nand4_1
X_06832_ _06145_ _06146_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__nor2_1
X_09551_ _02463_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__xor2_4
X_06763_ _05696_ _05707_ _05718_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__a21oi_1
X_08502_ _01395_ _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06694_ _03139_ _04972_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09482_ net283 _02401_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__or2_1
X_08433_ _01330_ _01331_ _01332_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08364_ net130 net131 net127 VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07315_ _00208_ _00217_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08295_ _01194_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07246_ _06339_ _06340_ _00147_ _00148_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07177_ net226 _03260_ _04752_ _00080_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09818_ _05498_ _01443_ _02064_ _03579_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__a22oi_1
X_09749_ _05969_ _02694_ _02695_ _03864_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a22oi_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _05913_ _05910_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or2b_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _04403_ _04420_ _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_84_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _05920_ _05921_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__and2_1
X_11642_ _04330_ _04331_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__and2b_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 data_in[115] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
X_11573_ _04136_ _04210_ _04697_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a21boi_4
Xinput29 data_in[125] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10524_ _02907_ _02916_ _02915_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__a21bo_1
X_10455_ _03467_ _03468_ _03470_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10386_ _06347_ _00879_ _02768_ _02766_ _02765_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__a32o_1
X_12125_ _05296_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nor2_1
X_12056_ _04827_ _05214_ _05225_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ _04074_ _04075_ _04064_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11909_ _05064_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__nand2_2
X_12889_ clknet_1_0__leaf_clk _00013_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07100_ _06412_ _06413_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08080_ _00976_ _00981_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07031_ net51 net60 net52 net61 VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08982_ _01871_ _01880_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__nand3_1
X_07933_ _02492_ _03864_ _00834_ net240 VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__nand4_1
X_07864_ _06077_ _06304_ _00763_ _00764_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__nand4_2
X_09603_ _02520_ _02533_ _02534_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__or3_1
X_06815_ net168 VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07795_ _00695_ _00696_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06746_ net68 _05520_ _05542_ _05509_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09534_ _01184_ _01790_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__or2_1
X_06677_ _04774_ _04785_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09465_ _01973_ _02382_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__nand3_1
X_08416_ _06077_ net213 net214 _03941_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__a22oi_2
X_09396_ _02307_ _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__xnor2_1
X_08347_ _00676_ _00685_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ _00243_ _00712_ _00714_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07229_ _00095_ _00131_ _00132_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__or3_4
XFILLER_0_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10240_ _03228_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10171_ _03131_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12812_ _06019_ _06024_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12743_ _05897_ _05898_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12674_ _05901_ _05902_ _05903_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11625_ _04738_ _04739_ _04751_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__or3_1
X_11556_ _01068_ _01629_ _04678_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10507_ _03526_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__xor2_2
XFILLER_0_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11487_ _04138_ _04164_ _04162_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10438_ _02832_ _02835_ _02834_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a21bo_1
X_10369_ _03364_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__xor2_2
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _05281_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__xor2_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _04357_ _04820_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06600_ _03941_ _02448_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and2_2
X_07580_ _03337_ net182 _00058_ _00481_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__nand4_1
X_06531_ net42 VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09250_ _01497_ _01504_ _01503_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08201_ _01019_ _01020_ _01101_ _01102_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__nor4_1
XFILLER_0_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06462_ _02415_ _02426_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__and2_1
X_09181_ _01436_ _01438_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08132_ net222 VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08063_ _00463_ _00964_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07014_ _06326_ _06327_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__and2_2
XFILLER_0_71_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput208 data_in[56] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
X_08965_ _01255_ _01258_ _01256_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__a21bo_1
Xinput219 data_in[66] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_2
X_07916_ _00816_ _00817_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__nand2_1
X_08896_ _01774_ _01224_ _01794_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__nand3_1
X_07847_ net153 VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_4
X_07778_ _06151_ _06274_ _00678_ _00679_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09517_ _04227_ net173 VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__and2_1
X_06729_ _05323_ _05334_ _05345_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__a21oi_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _02363_ _02364_ _01682_ _01684_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_109_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _01619_ _02288_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12390_ _05303_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__xnor2_1
X_11410_ _04499_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11341_ _00834_ _01385_ _01367_ _01987_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11272_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__or2_2
XFILLER_0_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10223_ _06274_ _00665_ _02551_ _02552_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__and4_1
X_10154_ _02485_ _02494_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__and2b_1
X_10085_ _01132_ _01133_ _01718_ _02398_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__a41o_4
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10987_ _04046_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__xor2_4
XFILLER_0_57_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12726_ _05790_ _05793_ _05959_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12657_ _05883_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11608_ _04265_ _04287_ _04285_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__a21o_2
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _05807_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11539_ _04658_ _04660_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _02800_ _01072_ _01075_ _01074_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__a31o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ _01007_ _01008_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__and2b_1
X_07701_ _00602_ net313 _00603_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__a21o_1
X_07632_ net36 _00533_ _00534_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09302_ net176 _00479_ _02203_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__a22o_1
X_07563_ _00452_ _00465_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__nand2_1
X_07494_ net63 VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__clkbuf_4
X_06514_ _02437_ _02987_ _02998_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__nand3_2
X_06445_ net85 VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__clkbuf_4
X_09233_ net105 net118 net119 net104 VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09164_ net84 VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08115_ _01001_ _01016_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09095_ _01366_ _01992_ _01993_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08046_ _00946_ _00947_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ net33 net227 net49 net225 VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__and4_2
XFILLER_0_99_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08948_ _01846_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__and2_1
X_08879_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__inv_2
X_10910_ _03962_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11890_ _04639_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10841_ _03290_ _03296_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10772_ _03816_ _03817_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12511_ _05489_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__xnor2_2
X_12442_ _05086_ _05087_ _05417_ _05418_ _05414_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12373_ _05566_ _05573_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11324_ _04384_ _04423_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__xor2_2
XFILLER_0_105_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11255_ _03829_ _03834_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__o21ai_4
X_10206_ _02555_ _03189_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__o21a_1
X_11186_ _04269_ _04271_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__and3_1
X_10137_ _03090_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__xnor2_4
X_10068_ _03045_ _03046_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12709_ _05857_ _05864_ _05862_ _05941_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09920_ _02851_ _02852_ _02882_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09851_ _02798_ _02806_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ _06086_ _06306_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__a21bo_1
X_09782_ _03732_ net66 _02731_ _03798_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a22oi_2
X_08802_ _01700_ _01701_ _01466_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__a21o_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _01630_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__xor2_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08664_ net182 net167 net197 _01563_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__and4_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ net218 net219 net229 VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08595_ _01494_ _01495_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__nor2_1
X_07546_ _00437_ _00448_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07477_ _00365_ _00378_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__and2_1
X_09216_ _06424_ _06410_ net72 _00421_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__nand4_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09147_ _02040_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09078_ _01547_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08029_ _00927_ _00928_ _00929_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11040_ _03533_ _03543_ _03542_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__a21bo_1
X_11942_ _04634_ _04695_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_87_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11873_ _04618_ _04629_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10824_ _03858_ _03873_ _03874_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10755_ _06134_ _01251_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10686_ _00270_ _01157_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12425_ _05362_ _05365_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a21oi_1
X_12356_ _05552_ _05554_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11307_ _04404_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__nor2_1
X_11238_ _04328_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__xor2_2
X_11169_ _03737_ _03700_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07400_ net199 net211 _06307_ _06306_ _06077_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ _01279_ _01280_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__xor2_2
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07331_ _06286_ _00233_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07262_ net257 VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkinv_4
X_07193_ net44 VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__buf_2
X_09001_ _01337_ _01339_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09903_ net100 net180 VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__and2_1
X_09834_ _02787_ _02788_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _02705_ _02711_ _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__nand3_1
X_06977_ _06288_ _06290_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__xnor2_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _02628_ _02636_ _02637_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__nand3_1
X_08716_ net224 VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08647_ _01545_ _01546_ _01468_ _01019_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a211oi_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ _01476_ _01477_ _00917_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__a21oi_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07529_ _03590_ net71 _00431_ _02657_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10540_ _02926_ _02938_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10471_ _02892_ _02900_ _02898_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _01629_ _02329_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12141_ _04944_ _04962_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__a21o_1
X_12072_ _01309_ _01288_ _02615_ _02592_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and4_1
X_11023_ _03551_ _03565_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a21o_2
X_11925_ _05081_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11856_ _00953_ _01563_ _01524_ _02215_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__nand4_1
X_10807_ _03320_ _03334_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11787_ _04929_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10738_ net98 net91 net99 net92 VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12408_ _05611_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__and2_1
X_10669_ _03132_ _03156_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12339_ _05192_ _05195_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__a21oi_2
X_06900_ _06205_ _06206_ _06213_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__o21ai_1
X_07880_ _00756_ _00311_ _00780_ _00781_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06831_ _06141_ _06144_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__and2_1
X_09550_ _02467_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__xnor2_2
X_06762_ _05696_ _05707_ _05718_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__and3_1
X_08501_ _00824_ _01401_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__xnor2_2
X_09481_ net283 _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and2_1
X_06693_ _04928_ _04961_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__xor2_4
X_08432_ _01330_ _01331_ _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08363_ net128 VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07314_ _00215_ _00216_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__nand2_1
X_08294_ _01180_ _00700_ _01193_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__and3_1
X_07245_ _06339_ _06340_ _00147_ _00148_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__nor4_1
XFILLER_0_131_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07176_ net220 VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09817_ _02769_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__xnor2_2
X_09748_ net242 VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _02616_ _02617_ _02614_ _01916_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__a211o_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _04417_ _04419_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__or2b_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12690_ _05858_ _05919_ _05869_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__or3_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _03774_ _04312_ _04770_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__o21ai_1
X_11572_ _04207_ _04209_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__or2b_1
Xinput19 data_in[116] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_4
XFILLER_0_107_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10523_ _03542_ _03543_ _03533_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10454_ net105 net120 VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__and2_1
X_10385_ _02758_ _02760_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12124_ _05299_ _05300_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__xnor2_1
X_12055_ _04827_ _05214_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a21oi_1
X_11006_ _04064_ _04074_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__nand3_1
X_11908_ _04193_ _04667_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12888_ clknet_1_0__leaf_clk _00012_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11839_ _00956_ _02132_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07030_ _02569_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08981_ _01877_ _01878_ _01879_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__nand3_1
X_07932_ net239 VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07863_ _06077_ net211 _00763_ _00764_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a22o_1
X_09602_ _02521_ _02532_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__and2_1
X_06814_ _06127_ _04259_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__a21bo_1
X_09533_ _01844_ _01846_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__nand2_2
X_07794_ _04435_ _00250_ _00693_ _00694_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__nand4_1
X_06745_ _05487_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06676_ _04752_ _03238_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__nand2_2
X_09464_ _02380_ _02381_ _01974_ _01975_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__a211o_1
X_08415_ _00775_ _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__xor2_2
X_09395_ _03084_ net48 VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08346_ _00215_ _00684_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08277_ _01177_ _00730_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__or2_1
X_07228_ _00127_ _00128_ _00130_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07159_ _03392_ _05191_ _05202_ _03381_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__a22o_1
X_10170_ _03132_ _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xor2_4
XFILLER_0_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12811_ _05999_ _05920_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__o21ai_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05898_ _05897_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _05901_ _05902_ _02185_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o21ai_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _04738_ _04739_ _04751_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11555_ _00530_ _01051_ _01653_ _02329_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11486_ _04121_ _04601_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o21ai_4
X_10506_ net176 net145 VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap308 _06269_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__buf_1
X_10437_ _02840_ _02841_ _02842_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10368_ _03365_ _03374_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _03297_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__xor2_1
X_12107_ _02694_ _01987_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__and3_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12038_ _04357_ _04820_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06530_ _02844_ _03172_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__xor2_4
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06461_ _02372_ _02405_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08200_ _01099_ _01100_ _00571_ _00573_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09180_ _02077_ _02078_ _02063_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08131_ _01024_ _01032_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08062_ _00952_ _00963_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__xor2_1
X_07013_ _06318_ _06325_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__nand2_1
Xinput209 data_in[57] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_4
X_08964_ _06152_ _00665_ _01861_ _01862_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__nand4_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07915_ _00807_ _00815_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__or2_1
X_08895_ _01774_ _01224_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a21o_1
X_07846_ _00744_ _00745_ _00746_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__a21oi_1
X_07777_ net130 net131 net126 _00677_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09516_ _02438_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__xor2_1
X_06728_ _05323_ _05334_ _05345_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__and3_1
X_09447_ _01682_ _01684_ _02363_ _02364_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__a211o_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06659_ _04216_ _04589_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__xnor2_1
X_09378_ _02286_ _02287_ _02282_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08329_ _06254_ net90 net91 _04413_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11340_ _01385_ _01367_ _01987_ _00834_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_120_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11271_ _04351_ _04364_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nor2_1
X_10222_ _06283_ _00210_ _00201_ _00677_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__and4_1
X_10153_ _02467_ _02476_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__o21ai_2
X_10084_ _03062_ _03063_ _02397_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10986_ _04052_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12725_ _05790_ _05793_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__o21ba_1
X_12656_ _05642_ _05709_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12587_ _05563_ _05576_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__a21oi_1
X_11607_ _04294_ _04433_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__a21o_2
XFILLER_0_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11538_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11469_ _04579_ _04580_ _04582_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _06224_ _00158_ _00159_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__and3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08680_ _01561_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__xnor2_2
X_07631_ net35 net43 net36 net42 VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__a22o_1
X_07562_ _00031_ _00464_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09301_ net174 net175 _00985_ net145 VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06513_ _02624_ _02965_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07493_ _00386_ _00395_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06444_ net94 VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09232_ net120 VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09163_ _01447_ _01452_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08114_ _01012_ _01015_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__xnor2_1
X_09094_ _01992_ _01993_ _01366_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08045_ _00423_ _00425_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09996_ _02304_ _02308_ _02305_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_110_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08947_ _01844_ _01845_ _01826_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__a21o_1
X_08878_ net166 net163 net164 net165 VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07829_ _00714_ _00715_ _00729_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__o21a_1
X_10840_ _03294_ _03295_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10771_ _06274_ _00210_ _01250_ net138 VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12510_ _05723_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__nor2_1
X_12441_ _05647_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12372_ _05567_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11323_ _04386_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11254_ _03830_ _03833_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10205_ _03190_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11185_ _03712_ _03714_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__or2_1
X_10136_ _03118_ _03119_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__nor2_2
X_10067_ _02197_ _02375_ _02374_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10969_ _04033_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__xor2_4
XFILLER_0_58_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12708_ _05601_ _05856_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12639_ _05623_ _05629_ _05627_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09850_ _02804_ _02805_ _02801_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__a21o_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ net209 net202 _06172_ net200 VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__a22o_1
X_09781_ net5 VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__clkbuf_4
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _01466_ _01700_ _01701_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__nand3_2
X_08732_ _00530_ _01631_ _01632_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__a21bo_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _02723_ _01562_ _01563_ net167 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_96_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ net217 _00516_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__nand2_1
X_08594_ _01485_ _01486_ _01493_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07545_ _00443_ _00444_ _00446_ _00447_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__a31o_1
X_07476_ _00365_ _00378_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ net80 net72 net81 net71 VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09146_ _02043_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09077_ _01429_ _01463_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08028_ _00927_ _00928_ _00929_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09979_ _02303_ _02323_ _02322_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o21bai_2
X_11941_ _04692_ _04694_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or2b_1
X_11872_ _04625_ _04627_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10823_ _03860_ _03284_ _03872_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10754_ _06253_ _01858_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10685_ _03720_ _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12424_ _05623_ _05629_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ _05552_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11306_ _00343_ net216 VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12286_ _05145_ _05146_ _05476_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11237_ _00200_ _03180_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__nand2_1
X_11168_ _03695_ _04232_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a21oi_2
X_10119_ _02466_ _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__xnor2_1
X_11099_ _04168_ _03628_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07330_ _00231_ _00232_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09000_ _01425_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__inv_2
X_07261_ _00162_ _00163_ _00164_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__a21oi_1
X_07192_ net33 net42 net35 net43 VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09902_ net111 net123 net177 net178 VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09833_ _02785_ _02786_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _02709_ _02710_ _02706_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__a21o_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _04358_ _06161_ _06289_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__o21a_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _02632_ _02633_ _02634_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a21o_1
X_08715_ _01606_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__xnor2_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _01468_ _01019_ _01545_ _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__o211a_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _00917_ _01476_ _01477_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__and3_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07528_ net72 VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07459_ _05914_ _03787_ _06373_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10470_ _02869_ _02871_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09129_ _03820_ _02481_ _00821_ _01397_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12140_ _04960_ _04946_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12071_ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11022_ _03562_ _03564_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__nor2_1
X_11924_ _01034_ _04123_ _05079_ _05080_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__nand4_1
XFILLER_0_87_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11855_ _01563_ _01524_ _02215_ _00953_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a22o_1
X_10806_ _03333_ _03321_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__and2b_1
X_11786_ _04475_ _04476_ _04477_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10737_ net91 _00703_ net92 _00238_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12407_ _05603_ _05610_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__nand2_1
X_10668_ _03113_ _03115_ _03112_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10599_ _03627_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12338_ _05534_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12269_ _05458_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__xor2_2
XFILLER_0_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06830_ _06141_ _06144_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__nor2_1
X_06761_ _02899_ _03502_ _03689_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__a21bo_1
X_06692_ _04939_ _03128_ _04950_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a21bo_1
X_08500_ _01396_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__xnor2_2
X_09480_ _02398_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__xor2_1
X_08431_ _00760_ _00768_ _00767_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08362_ _00682_ _00683_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07313_ _00212_ _00213_ _00214_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_73_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08293_ _01180_ _00700_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07244_ _00145_ _00146_ _05729_ _06341_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07175_ _04851_ _05049_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09816_ _06347_ _00879_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nand2_1
X_09747_ net241 VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__buf_2
X_06959_ _02229_ _04336_ _06157_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__and3_2
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _02614_ _01916_ _02616_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o211a_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _01527_ _01528_ _00955_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _03759_ _04313_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11571_ _04634_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10522_ _03533_ _03542_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10453_ _06437_ _00454_ net118 net119 VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand4_1
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10384_ _02796_ _02812_ _02810_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12123_ _04911_ _04913_ _04910_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__o21ba_1
X_12054_ _04824_ _05223_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11005_ _00059_ _03499_ _04071_ _04072_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__nand4_1
XFILLER_0_114_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11907_ _04662_ _04665_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__nand2_1
X_12887_ clknet_1_0__leaf_clk _00011_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dfxtp_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11838_ _04986_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__nand2_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11769_ _04910_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _01877_ _01878_ _01879_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__a21o_1
X_07931_ net244 net239 net240 net243 VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07862_ net209 _06172_ _06361_ net204 VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__nand4_2
X_09601_ _02521_ _02532_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nor2_1
X_06813_ _04227_ _04238_ _06127_ _02317_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__a22o_1
X_07793_ _04435_ net28 _00693_ _00694_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__a22o_1
X_09532_ _01775_ _01793_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a21o_2
X_06744_ _05487_ _05509_ net68 _05520_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__and4b_1
X_06675_ net217 _03238_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__and2_1
X_09463_ _01974_ _01975_ _02380_ _02381_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__o211ai_2
X_08414_ _01313_ _01314_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__or2b_1
X_09394_ _02304_ _02305_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08345_ _00323_ _00686_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08276_ _00728_ _00727_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__and2b_1
X_07227_ _00127_ _00128_ _00130_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__and3_4
XFILLER_0_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07158_ net176 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07089_ _06359_ _06360_ _06401_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12810_ _05999_ _05920_ _05998_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _05975_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ net263 _05734_ _05745_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _04749_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11554_ _04676_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11485_ _04130_ _04132_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__or2_1
X_10505_ net175 net156 VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10436_ _03434_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10367_ _03371_ _03373_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _02628_ _02637_ _02636_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__a21bo_1
X_12106_ _01385_ _01367_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nand2_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12037_ _05200_ _05205_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06460_ _02372_ _02405_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08130_ _01030_ _01031_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08061_ _00458_ _00962_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07012_ _06318_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08963_ _06152_ _00665_ _01861_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__a22o_1
X_07914_ _00807_ _00815_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _01775_ _01793_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__xnor2_1
X_07845_ _00744_ _00745_ _00746_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__and3_1
X_07776_ _04314_ _00210_ _00677_ _02218_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09515_ _01744_ _01746_ _01750_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06727_ _03326_ _03491_ _03304_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__o21ai_1
X_09446_ _02360_ _02362_ _02325_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__a21oi_2
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06658_ _04281_ _04578_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06589_ _03820_ _02470_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__nand2_1
X_09377_ _02282_ _02286_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__and3_1
X_08328_ _04424_ _06134_ _06284_ _00200_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08259_ _00175_ _00623_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11270_ _04351_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__and2_2
XFILLER_0_104_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10221_ _03211_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10152_ _02474_ _02475_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10083_ _01712_ net286 _02393_ _02395_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_97_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10985_ _03453_ _03460_ _03459_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__o21ba_2
X_12724_ _05771_ _05779_ _05778_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12655_ _05708_ _05705_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12586_ _05565_ _05574_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__and2b_1
X_11606_ _04432_ _04295_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__and2b_1
X_11537_ _00544_ _01072_ _01667_ _03019_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11468_ _04579_ _04580_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11399_ _04505_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__xnor2_2
X_10419_ _03317_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__xor2_4
XFILLER_0_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ net42 net35 net43 VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07561_ _00461_ _00462_ _00463_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09300_ net175 net134 net145 net174 VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__a22o_1
X_06512_ _02976_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__inv_2
X_07492_ _00393_ _00394_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06443_ net121 VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09231_ _02129_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09162_ _00917_ _01476_ _01477_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08113_ _01013_ _01014_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09093_ _01990_ _01991_ _01381_ _01383_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_71_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08044_ _00944_ _00945_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09995_ _02283_ _02287_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__nand2_1
X_08946_ _01826_ _01844_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__nand3_1
X_08877_ net162 VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_4
X_07828_ _00714_ _00715_ _00729_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__nor3_1
XFILLER_0_67_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07759_ _00224_ _00262_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10770_ _00210_ _01250_ _03210_ _06274_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ _02789_ _03106_ net223 net234 VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__nand4_1
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12440_ _05643_ _05401_ _05646_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__nor3_1
XFILLER_0_75_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12371_ _05569_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11322_ _04388_ _04421_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11253_ _04335_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__xor2_2
XFILLER_0_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10204_ _02546_ _03193_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__xor2_1
X_11184_ _00617_ _02464_ _03709_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand3_1
X_10135_ _03091_ _03092_ _03116_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__and3_1
X_10066_ _02890_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10968_ _03439_ _03441_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__and2_2
X_12707_ _05800_ _05801_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__or2b_1
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10899_ _03954_ _03955_ _03956_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a21oi_1
X_12638_ _05857_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _05785_ _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _01697_ _01699_ _01105_ net291 VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06992_ net200 net209 _06172_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__and3_1
X_09780_ _02728_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__nand2_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _04906_ net46 net47 net33 VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a22o_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ net145 VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07613_ net230 VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_4
X_08593_ _01485_ _01486_ _01493_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07544_ _00443_ _00444_ _00446_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07475_ _06371_ _00377_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09214_ _01471_ _01473_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09145_ _02470_ _00850_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09076_ _01462_ _01460_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08027_ _00445_ _00444_ _00443_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09978_ _02290_ _02291_ _02292_ _02296_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__a31o_2
X_08929_ net25 net21 VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__and2_1
X_11940_ _05053_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11871_ _04975_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__xor2_2
X_10822_ _03860_ _03284_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10753_ _03213_ _03223_ _03222_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_94_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10684_ _03707_ _03708_ _03719_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__or3b_1
X_12423_ _05627_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__nor2_1
X_12354_ _04824_ _05223_ _05221_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11305_ _03885_ _03888_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12285_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11236_ _04326_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__xnor2_2
X_11167_ _04229_ _04231_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__nor2_1
X_10118_ _03098_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__xor2_1
X_11098_ _04174_ _04176_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__xnor2_1
X_10049_ _03018_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07260_ net278 _06218_ _06222_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__a21bo_1
X_07191_ _00093_ _00094_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09901_ net123 net177 net178 net111 VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09832_ _02785_ _02786_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__nor2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _02706_ _02709_ _02710_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__nand3_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _01613_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__and2b_1
X_06975_ _02240_ _06159_ _06158_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__nand3_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _02632_ _02633_ _02634_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__nand3_1
Xrebuffer10 _00584_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _01515_ _01516_ _01543_ _01544_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _01474_ _01475_ _01469_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__a21o_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07527_ _00428_ _00429_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__or2_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07458_ _00354_ _00360_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07389_ _02383_ _04139_ _06311_ _00291_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__nand4_2
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09128_ _02026_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09059_ _01901_ _01957_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__nor3_2
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12070_ _01288_ _02615_ _02592_ _01309_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11021_ _04023_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11923_ _01034_ _04123_ _05079_ _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11854_ _04100_ _04616_ _05004_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__o21ai_2
X_10805_ _03277_ _03302_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11785_ _03966_ _04480_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10736_ _06159_ _03180_ _03179_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10667_ _03158_ _03246_ _03245_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_36_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12406_ _05603_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ _03620_ _03626_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12337_ _05522_ _05533_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12268_ _05024_ _05103_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11219_ _00239_ _00706_ _00647_ _01181_ _03756_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a41o_1
X_12199_ _05003_ _05017_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput190 data_in[3] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
X_06760_ _05356_ _05367_ _05685_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__o21ai_1
X_06691_ net112 net256 net179 net245 VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08430_ _01328_ _01329_ _01321_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08361_ _01254_ _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07312_ _00212_ _00213_ _00214_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__or3b_2
XFILLER_0_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08292_ _01185_ _01192_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07243_ _05729_ _06341_ _00145_ _00146_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__o211a_2
XFILLER_0_61_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07174_ _05016_ _05038_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09815_ _02765_ _02766_ _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__a21bo_1
X_09746_ _02691_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__xor2_4
X_06958_ _06260_ _06271_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__xnor2_1
X_09677_ _03941_ net216 _02615_ _04139_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__a22o_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _00955_ _01527_ _01528_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__or3_1
X_06889_ _06125_ _06126_ _06200_ _06202_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _01430_ _01459_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ _04692_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10521_ _03540_ _03541_ _03534_ _03536_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10452_ net107 net118 net119 net106 VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10383_ _03389_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__nand2_1
X_12122_ _05297_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__or2_1
X_12053_ _05221_ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nor2_1
X_11004_ _00059_ _03499_ _04071_ _04072_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__a22o_1
X_11906_ _05054_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12886_ clknet_1_0__leaf_clk _00010_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dfxtp_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11837_ _00910_ _01520_ _01484_ _02164_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__nand4_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _01410_ _01397_ _02731_ _00821_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10719_ _03755_ _03756_ _03757_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11699_ _04814_ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__xnor2_2
Xrebuffer1 _00581_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07930_ _00829_ _00831_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07861_ _06172_ _06361_ net204 net209 VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09600_ _02522_ _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__xor2_1
X_07792_ _06138_ net26 net18 _06264_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06812_ net159 VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__buf_2
X_06743_ net79 VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09531_ _01776_ _01792_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06674_ _03227_ _03260_ _04752_ _02855_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__a22o_1
X_09462_ _02378_ _02379_ _02109_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__a21o_1
X_08413_ _01310_ _01312_ _00759_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__a21o_1
X_09393_ _04906_ net36 net46 net47 VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08344_ _01243_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08275_ _00278_ _00654_ _01175_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__o21ai_2
X_07226_ _04895_ _05005_ _00129_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07157_ _02723_ _02734_ _00058_ _00059_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07088_ _06359_ _06360_ _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__or3_4
XFILLER_0_30_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09729_ _05980_ net249 _02005_ _02004_ _00834_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _05973_ _05974_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ net264 _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__xor2_2
XFILLER_0_96_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _01777_ _01754_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11553_ _01051_ _01653_ net40 _00530_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11484_ _04130_ _04132_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__and2_1
X_10504_ _02895_ _02897_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__or2b_2
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10435_ _03446_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10366_ _05750_ _02733_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12105_ _01367_ _02695_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__nand2_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _03290_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12036_ _05203_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__xor2_4
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12869_ _06100_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__nor2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08060_ _00476_ _00961_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07011_ _06323_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08962_ net125 net133 net126 net135 VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__nand4_1
X_07913_ _00808_ _00814_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__xnor2_1
X_08893_ _01776_ _01792_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__xnor2_1
X_07844_ _00316_ _00317_ _00315_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07775_ net127 VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__buf_2
X_09514_ _02435_ _02436_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__nand2_1
X_06726_ _05071_ _05312_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__nand2_1
X_09445_ _02325_ _02360_ _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__and3_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06657_ _04556_ _04567_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__or2_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06588_ net253 VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__clkbuf_4
X_09376_ net227 net224 _02283_ _02285_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nand4_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08327_ _00203_ _00668_ _00669_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08258_ _01156_ _01158_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__xnor2_1
X_07209_ net256 net179 net190 net245 VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08189_ _01071_ _01089_ _01090_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nor3_1
X_10220_ _06152_ _06274_ _01250_ _03210_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__and4_2
XFILLER_0_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10151_ _02511_ _02513_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nand2_2
Xoutput280 net280 VGND VGND VPWR VPWR data_out[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10082_ net286 _01715_ _01717_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10984_ _04049_ _04050_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12723_ _05768_ _05814_ _05956_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12654_ _05852_ _05881_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12585_ _05798_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11605_ _04263_ _04289_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__or2b_1
XFILLER_0_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11536_ _01072_ _01667_ _03019_ _00544_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11467_ _00062_ _02215_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11398_ _03990_ _03992_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__nand2_1
X_10418_ _03428_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10349_ _03351_ _03352_ _02727_ _02729_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _01181_ _02498_ _01784_ _01217_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ _00067_ _00460_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06511_ _02624_ _02965_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nor2_1
X_07491_ net59 _00387_ _00391_ _00392_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__a22o_1
X_09230_ _05520_ _01487_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nand2_1
X_06442_ net130 VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09161_ _01442_ _01454_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09092_ _01381_ _01383_ _01990_ _01991_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08112_ _00497_ _00496_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08043_ _00943_ _00941_ _00942_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09994_ _02955_ _02964_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__xor2_2
X_08945_ _01827_ _01828_ _01843_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08876_ _00709_ _01206_ _01208_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__o21ba_1
X_07827_ _00727_ _00728_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__xor2_1
X_07758_ _00196_ _00223_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06709_ _02723_ _05093_ _05104_ _05126_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__nand4_2
X_07689_ _00589_ _00590_ _00147_ net322 VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09428_ net12 _01666_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09359_ net219 net231 net232 net218 VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a22oi_2
X_12370_ _05570_ _03859_ _05253_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__mux2_4
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11321_ _04403_ _04420_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11252_ _04343_ _04344_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _03191_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__xor2_1
X_11183_ _00617_ _01188_ _02464_ _00171_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a22o_1
X_10134_ _03091_ _03092_ _03116_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__a21oi_1
X_10065_ _03041_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__xor2_4
XFILLER_0_106_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10967_ _04031_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__xor2_4
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10898_ _03954_ _03955_ _03956_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12706_ _05798_ _05806_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__nand2_1
X_12637_ _05862_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12568_ _05251_ _05786_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11519_ _01034_ _01023_ _01617_ _01603_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__and4_1
X_12499_ _05710_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _02459_ _06304_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ net33 _04906_ net47 VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__and3_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ net197 VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__buf_2
X_07612_ _00512_ _00514_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08592_ _01491_ _01492_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07543_ _00445_ _06419_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07474_ _00369_ _00376_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _01474_ _01476_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09144_ _03798_ net4 VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09075_ _01466_ _01700_ _01701_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and3_1
X_08026_ _00925_ _00926_ _00920_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09977_ _02945_ _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__nor2_2
X_08928_ _01216_ _01219_ _01220_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08859_ _01735_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11870_ _04977_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__xor2_2
X_10821_ _03866_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10752_ _03190_ _03195_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10683_ _03707_ _03708_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__o21bai_1
X_12422_ _04539_ _05353_ _05626_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12353_ _05550_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11304_ _04400_ _04401_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12284_ _05145_ _05146_ _05476_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11235_ _03780_ _03783_ _03781_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11166_ _04236_ _04241_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a21oi_1
X_11097_ _00097_ _02329_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__and3_1
X_10117_ _00270_ net171 VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nand2_1
X_10048_ _03023_ _03024_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11999_ _01188_ _01754_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07190_ _04818_ _00092_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09900_ net89 _01524_ _02170_ _02171_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09831_ _02059_ _02098_ _02097_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _03820_ _02019_ _02707_ _02708_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nand4_2
X_06974_ _06282_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _01611_ _01612_ _01607_ _01608_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__a211o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _01920_ _01922_ _01921_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08644_ _01515_ _01516_ _01543_ _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__nand4_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _01469_ _01474_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__nand3_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07526_ _06412_ _00427_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__nor2_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07457_ _00356_ _00358_ _00359_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07388_ net143 VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09127_ _02024_ _02025_ _02022_ _02023_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09058_ _01955_ _01956_ _01902_ _01376_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08009_ _02646_ _00910_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11020_ _04089_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__or2b_2
Xmax_cap290 _01111_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11922_ _01023_ _01617_ _01603_ _03580_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__nand4_2
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _04109_ _04111_ _04614_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__a21o_1
X_10804_ _03301_ _03300_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11784_ _04926_ _04927_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10735_ _03177_ _03178_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10666_ _03118_ _03701_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__or2_2
X_12405_ _05607_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10597_ _03620_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12336_ _05522_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12267_ _05100_ _05102_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__nor2_1
X_11218_ _04306_ _01784_ _00239_ _04304_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__and4b_1
X_12198_ _05015_ _05006_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__or2b_1
X_11149_ _03695_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput180 data_in[30] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_2
Xinput191 data_in[40] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
X_06690_ net179 VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08360_ _01259_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07311_ _06276_ _06278_ _06275_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08291_ _01190_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07242_ _06406_ _06407_ _00143_ _00144_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07173_ _00075_ _00076_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09814_ net61 net57 net58 net60 VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__a22o_1
X_09745_ _06384_ _00830_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__nand2_2
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06957_ net308 _06270_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__nor2_1
X_09676_ _03941_ _04139_ net216 _02615_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nand4_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06888_ _06125_ _06126_ _06200_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__nor4_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ net78 net180 _01525_ _01526_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__and4_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _01431_ _01458_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__xor2_2
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08489_ _01387_ _01388_ _01389_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__a21o_1
X_07509_ _00383_ _00384_ _00411_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10520_ _03534_ _03536_ _03540_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10451_ _05520_ _02799_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10382_ _02764_ _02780_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12121_ _01410_ _01397_ _02731_ _02019_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__and4_1
X_12052_ _05215_ _04861_ _05220_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__nor3_1
X_11003_ _04068_ _04069_ _04070_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a21o_1
X_11905_ _05055_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__xnor2_4
X_12885_ clknet_1_0__leaf_clk _00009_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dfxtp_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11836_ _01520_ _01484_ _02164_ _00910_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _00821_ _01410_ _01397_ _02731_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10718_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_125_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11698_ _04831_ _04833_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__xor2_2
XFILLER_0_113_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer2 _01688_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
X_10649_ _03075_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12319_ _05493_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_1
X_07860_ net200 net211 _00299_ _00300_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__and4_1
X_07791_ net26 net18 net27 net17 VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a22o_1
X_06811_ _06122_ _06123_ _06124_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a21oi_1
X_09530_ _01817_ _01849_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__or2_2
X_06742_ _03579_ _03590_ _05498_ _02657_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__a22o_1
X_09461_ _02109_ _02378_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__nand3_1
X_06673_ net219 VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__clkbuf_4
X_08412_ _00759_ _01310_ _01312_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__and3_1
X_09392_ net36 _00530_ _01051_ _04906_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08343_ _01226_ _01242_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08274_ _00256_ _00653_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07225_ _03150_ _04994_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07156_ _02723_ _00058_ _00059_ _02734_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07087_ _06399_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__or2_2
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09728_ _01989_ _01991_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__or2_1
X_07989_ _00428_ _00889_ _00890_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__nand3_1
X_09659_ _06171_ _06319_ _00774_ net146 VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nand4_1
XFILLER_0_97_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05747_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11621_ _04746_ _04748_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11552_ _03624_ _04196_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10503_ _02948_ _02978_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11483_ _04532_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10434_ _03444_ _03445_ _03435_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a21o_1
X_10365_ _05750_ net66 _02733_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12104_ _04443_ _04899_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _03294_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12035_ _01251_ _03180_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12868_ net319 _06103_ _06107_ _06100_ _02185_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11819_ _04493_ _04521_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _06038_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07010_ _06321_ _06322_ _06181_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08961_ net133 net126 net135 net125 VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a22o_1
X_07912_ _00809_ _00813_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__xnor2_1
X_08892_ _01783_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__xnor2_1
X_07843_ net140 net152 _00742_ _00743_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__nand4_1
X_07774_ _00674_ _00675_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09513_ _02433_ _02434_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__nand2_1
X_06725_ _05071_ _05312_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__or2_1
X_09444_ _02358_ _02359_ _02326_ _01680_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__a211o_2
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06656_ _02295_ _04545_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and2_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06587_ _03798_ _02481_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__nand2_1
X_09375_ net227 net224 _02283_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08326_ _00721_ _00722_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08257_ _02328_ _01157_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07208_ net245 net256 net179 net190 VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__nand4_1
X_08188_ _01086_ _01087_ _01088_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07139_ _00041_ _00042_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10150_ _03133_ _03134_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__nand2_4
Xoutput270 net270 VGND VGND VPWR VPWR data_out[20] sky130_fd_sc_hd__clkbuf_4
Xoutput281 net281 VGND VGND VPWR VPWR data_out[5] sky130_fd_sc_hd__clkbuf_4
X_10081_ _03059_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__nor2_1
X_10983_ _03455_ _03457_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__and2_2
X_12722_ _05813_ _05770_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12653_ _05853_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12584_ _05803_ _05804_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11604_ _04288_ _04264_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11535_ _04636_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11466_ _05202_ _01563_ _03532_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11397_ _04503_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__xor2_2
X_10417_ _03318_ _03427_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nor2_1
X_10348_ _02727_ _02729_ _03351_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a211o_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _03255_ _03276_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__xnor2_2
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _04310_ _04786_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07490_ _02569_ _00387_ _00391_ _00392_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__nand4_2
XFILLER_0_75_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06510_ _02943_ _02954_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__or2_1
X_06441_ net15 VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09160_ _00885_ _01453_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09091_ _01988_ _01989_ net208 _01986_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08111_ _00494_ _00495_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08042_ _00941_ _00942_ _00943_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _02962_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ _01827_ _01828_ _01843_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08875_ _01185_ _01192_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__and2_1
X_07826_ _06286_ _00233_ _00235_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__o21a_1
X_07757_ _00657_ _00658_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06708_ _02723_ _05093_ _05104_ _05126_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07688_ _00147_ net288 _00589_ _00590_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__o211ai_4
X_09427_ _02341_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__xnor2_1
X_06639_ _02273_ _04358_ _04369_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__and3_1
X_09358_ _01642_ _01643_ _01069_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__or3b_1
XFILLER_0_136_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08309_ _01208_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__or2_1
X_11320_ _04417_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09289_ _02157_ _02158_ _02188_ _02189_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11251_ _04342_ _04337_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__or2b_1
X_10202_ net97 net92 VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__nand2_1
X_11182_ _03723_ _03724_ _03720_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__o21a_1
X_10133_ _03114_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10064_ _02264_ _02370_ _02369_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_89_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10966_ _01487_ _00937_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10897_ _03346_ _03354_ _03353_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12705_ _05775_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__xor2_4
XFILLER_0_122_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12636_ _05607_ _05611_ _05861_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12567_ _05251_ _05568_ _05786_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11518_ _01023_ _01617_ _01603_ _01034_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12498_ _05349_ _05461_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__a21oi_1
X_11449_ _04053_ _04052_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__or2b_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ net211 VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__buf_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _01559_ _01560_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__or2_1
X_07611_ _04785_ _00081_ _00513_ _00510_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__or4_1
X_08591_ _05520_ _00431_ _01489_ _01490_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__nand4_2
X_07542_ _03524_ _02646_ _05444_ _06416_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07473_ _00374_ _00375_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09212_ _01552_ _01596_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09143_ _02041_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09074_ _01700_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08025_ _00920_ _00925_ _00926_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09976_ _02255_ _02257_ _02944_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__and3_1
X_08927_ _00705_ _01215_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08858_ _01756_ _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07809_ _00704_ _00705_ _00707_ _00709_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a22oi_1
X_08789_ _01046_ _01098_ _01097_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__o21bai_1
X_10820_ _03869_ _03870_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10751_ _02546_ _03193_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10682_ _03717_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand2_1
X_12421_ _04539_ _05353_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12352_ _05218_ _05549_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11303_ _04399_ _04398_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12283_ _05148_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11234_ _04323_ _04324_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11165_ _04233_ _04235_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__nor2_1
X_11096_ _04862_ _01653_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__nand2_1
X_10116_ _03096_ _03097_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
X_10047_ _02344_ _02346_ _02345_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11998_ _05157_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__xnor2_1
X_10949_ _03982_ _04012_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12619_ _05842_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09830_ _02750_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__xnor2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _03820_ net14 _02707_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a22o_1
X_06973_ _06285_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__and2_2
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _01607_ _01608_ _01611_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__o211a_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _02629_ _02630_ _02631_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__nand3_1
XFILLER_0_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08643_ _01539_ _01540_ _01542_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _01472_ _01473_ _00913_ _00915_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _06412_ _00427_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__and2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07456_ _06373_ _00355_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07387_ _06310_ _06316_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09126_ _02022_ _02023_ _02024_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _01902_ _01376_ _01955_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08008_ net118 VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap291 _01107_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_2
X_09959_ _02276_ _02277_ _01610_ _01611_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11921_ _01617_ _01603_ _03580_ _01023_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a22o_1
X_11852_ _04583_ _04585_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__nand2_1
X_10803_ _03335_ _03384_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11783_ _04476_ _04925_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10734_ _03774_ _03775_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10665_ _03090_ _03120_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12404_ _05604_ _05606_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10596_ _03621_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12335_ _05530_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12266_ _05388_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11217_ _00239_ _01784_ _04305_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__o2bb2a_1
X_12197_ _05380_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__and2_1
X_11148_ _04229_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__xor2_2
Xinput170 data_in[252] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
Xinput181 data_in[31] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
X_11079_ _04153_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__xor2_1
Xinput192 data_in[41] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07310_ net124 net132 _00209_ _00211_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08290_ _01189_ _00270_ net168 _01186_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__and4b_1
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07241_ _06406_ _06407_ _00143_ _00144_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__nand4_2
XFILLER_0_116_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07172_ _00046_ _00074_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09813_ net60 net61 net57 VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09744_ _01385_ _02688_ _02689_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__a21bo_1
X_06956_ _06262_ _06263_ _06267_ _06268_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__o22a_1
X_09675_ net147 VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__clkbuf_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06887_ _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__inv_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _02745_ _01524_ _01525_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__a22oi_2
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _01432_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__xnor2_2
X_08488_ net246 _00834_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07508_ _00408_ _00410_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07439_ _06389_ _06390_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10450_ _03461_ _03462_ _03463_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09109_ net244 net241 net242 _02492_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10381_ _02779_ _02777_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _01397_ _02731_ _02019_ _01410_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12051_ _05215_ _04861_ _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11002_ _04068_ _04069_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__nand3_1
X_11904_ _04664_ _05059_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__xor2_4
XFILLER_0_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12884_ clknet_1_0__leaf_clk _00008_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11835_ _04982_ _04984_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__nand2_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _00830_ _02695_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10717_ _03755_ _03756_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__or3b_1
XFILLER_0_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11697_ _04349_ _04368_ _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 _01688_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_1
XFILLER_0_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10648_ _03681_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10579_ _00107_ _01629_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12318_ _05495_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__xnor2_4
X_12249_ _04606_ _05434_ _05437_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__nor3_1
X_07790_ _00690_ _00691_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__nor2_2
X_06810_ _06122_ _06123_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__and3_1
X_06741_ net70 VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09460_ _02376_ _02377_ _01695_ _02110_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__a211o_1
X_08411_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__inv_2
X_06672_ net228 VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__buf_2
X_09391_ _01634_ _01641_ _01640_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08342_ _01226_ _01242_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08273_ _00795_ _00797_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__nand2_1
X_07224_ _00125_ _00126_ _00105_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07155_ net111 VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07086_ _06366_ _06398_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07988_ _00887_ _00888_ _00878_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a21o_1
X_09727_ _02008_ _02016_ _02015_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__o21bai_2
X_06939_ net97 VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09658_ net151 _00774_ net146 net150 VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _01253_ _01812_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__a21oi_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _01496_ _01508_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__nand3_4
XFILLER_0_77_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _01777_ _01157_ _04276_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__a31o_1
X_11551_ _04191_ _04195_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10502_ _02977_ _02949_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11482_ _04596_ _04597_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10433_ _03435_ _03444_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__and3_1
X_10364_ _03368_ _03369_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12103_ _04458_ _04898_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__nand2_1
X_10295_ _02629_ _02631_ _02630_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__a21bo_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12034_ _01835_ _01858_ _05201_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__and3_2
XFILLER_0_125_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12867_ net274 net275 VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nand2_1
X_11818_ _04520_ _04495_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__and2b_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _06035_ _06037_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11749_ _04522_ _04525_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08960_ _01857_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07911_ _00811_ _00812_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__nand2_1
X_08891_ _01184_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__xnor2_2
X_07842_ net140 net152 _00742_ _00743_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07773_ _00670_ _00671_ _00673_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o21ai_1
X_09512_ _02433_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__or2_1
X_06724_ _05290_ _05301_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__or2_1
X_09443_ _02326_ _01680_ _02358_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__o211ai_2
X_06655_ _02295_ _04545_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__nor2_1
X_09374_ net32 net49 net225 net226 VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__a22o_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06586_ net7 VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08325_ _01224_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08256_ net172 VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__buf_2
X_07207_ net112 net12 VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08187_ _01086_ _01087_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07138_ _05597_ _00040_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__or2_1
X_07069_ net247 VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput260 net260 VGND VGND VPWR VPWR data_out[11] sky130_fd_sc_hd__clkbuf_4
Xoutput271 net271 VGND VGND VPWR VPWR data_out[21] sky130_fd_sc_hd__clkbuf_4
Xoutput282 net282 VGND VGND VPWR VPWR data_out[6] sky130_fd_sc_hd__clkbuf_4
X_10080_ _02391_ _02393_ _03058_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10982_ _04047_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12721_ _05756_ _05759_ _05762_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a21o_2
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12652_ _05878_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11603_ _04261_ _04290_ _04728_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12583_ _05799_ _05616_ _05802_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11534_ _04653_ _04654_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11465_ _00479_ _03499_ _04576_ _04577_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__nand4_1
X_10416_ _03318_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11396_ _00879_ _01434_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10347_ _03347_ _03349_ _03350_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _03274_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _04806_ _04810_ _04812_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap1 _01115_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_2
XFILLER_0_119_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06440_ net24 VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__clkbuf_4
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09090_ net208 _01986_ _01988_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__o2bb2a_1
X_08110_ _01010_ _01011_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08041_ _00433_ _00435_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09992_ _02960_ _02961_ _02956_ _02277_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__a211o_1
X_08943_ _01834_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08874_ _00710_ _01222_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__nand2_1
X_07825_ _00716_ _00726_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__xor2_2
X_07756_ _00639_ _00640_ _00656_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__or3_1
X_06707_ _03337_ _02712_ _03348_ _05115_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__nand4_4
X_09426_ _04939_ _01072_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nand2_1
X_07687_ _00339_ _00340_ _00587_ _00588_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06638_ _04292_ _02240_ _04325_ _04347_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__a22o_1
X_09357_ _00513_ _01036_ _01622_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06569_ _03579_ _02657_ _03590_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _02157_ _02158_ _02188_ _02189_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__and4_1
X_08308_ _00694_ _00696_ _01207_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08239_ _00734_ _00736_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11250_ _04337_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10201_ _06254_ net93 VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__nand2_1
X_11181_ _03744_ _03767_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__or2b_1
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10132_ _06127_ net173 VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__nand2_1
X_10063_ _02947_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12704_ _05251_ _05786_ _05787_ _05785_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__a2bb2o_2
X_10965_ net75 _04028_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a21bo_1
X_10896_ _03951_ _03953_ _03945_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12635_ _05607_ _05611_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12566_ _01872_ _03210_ _05244_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11517_ _04167_ _04179_ _04178_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12497_ _05458_ _05460_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11448_ _04555_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__xnor2_4
X_11379_ _04481_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07610_ net226 _03260_ _00080_ _00507_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__and4_1
X_08590_ _05520_ _00431_ _01489_ _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a22o_1
X_07541_ _00441_ _00442_ _00030_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07472_ _03853_ _05969_ _06386_ _06385_ _06384_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09211_ _01543_ _01545_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__nand2_1
X_09142_ net50 net6 net66 net5 VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09073_ _01971_ _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08024_ _00923_ _00924_ _00456_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09975_ _02255_ _02257_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__a21oi_2
X_08926_ _01819_ _01825_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08857_ _01753_ _01755_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07808_ _00704_ _00705_ _00707_ _00709_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__and4_1
X_08788_ _01626_ _01627_ _01686_ _01687_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07739_ _06265_ _00254_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__nor2_1
X_10750_ _03777_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09409_ _02320_ _02321_ _01657_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10681_ _03715_ _03716_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12420_ _02799_ _04953_ _05625_ _02064_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12351_ _05218_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11302_ _04398_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__and2b_1
X_12282_ _05473_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11233_ _00672_ _01835_ _04320_ _04322_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a22oi_1
X_11164_ _04248_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
X_11095_ _04171_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__xor2_1
X_10115_ net169 _00171_ _01777_ _01188_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand4_1
X_10046_ _03021_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__nor2_2
X_11997_ _05160_ _05161_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10948_ _03983_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10879_ _03921_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__xor2_4
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12618_ _05694_ _05840_ _05841_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12549_ _05562_ _05580_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09760_ net254 _06375_ net11 net13 VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__nand4_2
X_06972_ _02229_ _02240_ _06283_ _06284_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__nand4_4
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _02629_ _02630_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__a21o_1
X_08711_ _04752_ _00516_ _01609_ _01610_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a22o_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08642_ _01539_ _01540_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__nand3_2
XFILLER_0_83_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08573_ _00913_ _00915_ _01472_ _01473_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ _00425_ _00426_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__nor2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07455_ _03798_ net255 _00357_ _02470_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07386_ _06182_ _06317_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09125_ _05914_ _00822_ _01406_ _01407_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09056_ _01934_ _01935_ _01954_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_102_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08007_ _00093_ _00500_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap292 _00736_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_1
X_09958_ _02244_ _02246_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_2
X_08909_ _04424_ _06134_ _00672_ net92 VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__nand4_1
X_09889_ _02846_ _02847_ _02815_ _02153_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__a211o_1
X_11920_ _04673_ _04683_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11851_ _04568_ _04588_ _04587_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__o21ba_1
X_10802_ _03380_ _03383_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__or2_1
X_11782_ _04476_ _04925_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10733_ _03163_ _03770_ _03773_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10664_ _03126_ _03314_ _03698_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21o_2
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10595_ _03622_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12403_ _05604_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12334_ _04781_ _05189_ _05529_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12265_ _05453_ _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__xnor2_2
X_11216_ _00706_ _00647_ _01217_ _01181_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__and4_1
X_12196_ _05369_ _05379_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11147_ _03125_ _03674_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput171 data_in[253] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xinput160 data_in[243] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
X_11078_ _00107_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand2_1
Xinput182 data_in[32] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
Xinput193 data_in[42] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
X_10029_ _04939_ net45 _02340_ _02338_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07240_ _00141_ _00142_ _06408_ _05696_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07171_ _00046_ _00074_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09812_ net58 VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__clkbuf_4
X_09743_ net239 net248 net240 net247 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06955_ _06262_ _06263_ _06267_ _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__nor4_1
X_09674_ _06086_ _06362_ _00297_ _00757_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__and4_1
X_06886_ _06199_ _06197_ _06198_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__nand3_2
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ net89 net100 net177 net178 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__nand4_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _01455_ _01456_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__xor2_2
XFILLER_0_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07507_ _00409_ _06359_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__nor2_1
X_08487_ _02492_ _03864_ net240 net241 VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__nand4_1
XFILLER_0_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07438_ _06409_ _00039_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07369_ _00271_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__inv_2
X_09108_ _02006_ _02007_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10380_ _02814_ _02850_ _02848_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09039_ net140 _06177_ net153 net154 VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12050_ _05218_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11001_ _03489_ _03492_ _03490_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11903_ _04660_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12883_ clknet_1_0__leaf_clk _00007_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dfxtp_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11834_ _04978_ _04981_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__or2_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11765_ _04905_ _04907_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11696_ _04367_ _04350_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__or2b_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _03144_ _03145_ _03143_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10647_ _03076_ _03077_ _03680_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer4 net325 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
X_10578_ _03604_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12317_ _05511_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__nand2_2
X_12248_ _04606_ _05434_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12179_ _04993_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2_1
X_06740_ net69 net76 net77 net70 VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06671_ _03216_ _03249_ _03271_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nand3_2
X_08410_ net148 net149 net144 net146 VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__and4_1
X_09390_ _02300_ _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08341_ _01240_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08272_ _01138_ _01172_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__xnor2_2
X_07223_ _00105_ _00125_ _00126_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__or3_4
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07154_ net194 VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07085_ _06366_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07987_ _00878_ _00887_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__nand3_1
X_09726_ _01992_ _01995_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__nand2_1
X_06938_ _06148_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09657_ _01944_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__inv_2
X_06869_ _06182_ _06183_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _01813_ _01807_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__and2b_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _01505_ _01506_ _01507_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__a21o_1
X_08539_ _01437_ _01438_ _01433_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _03610_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__or2_2
XFILLER_0_135_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10501_ _02925_ _02941_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11481_ _04594_ _04595_ _04533_ _04535_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10432_ _03442_ _03443_ _03437_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10363_ net10 _00850_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12102_ _04916_ _04918_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__and2b_1
X_10294_ _03291_ _03292_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nor2_1
X_12033_ _00703_ _01251_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12866_ _06106_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__clkbuf_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11817_ _04940_ _04964_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__xor2_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12797_ _06035_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11748_ _04764_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__xor2_4
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11679_ _04805_ _04811_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07910_ _02448_ _00810_ _00368_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__a21o_1
X_08890_ _01788_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__or2_2
X_07841_ _06177_ net150 net142 net151 VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__nand4_2
X_07772_ _00670_ _00671_ _00673_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__or3_2
XFILLER_0_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09511_ _06127_ _01157_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__and2_1
X_06723_ _03436_ _05279_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09442_ _02356_ _02357_ _02337_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__o21ai_2
X_06654_ _04523_ _04534_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__or2_1
X_06585_ net253 net6 net7 VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__and3_1
X_09373_ net32 net226 net49 net225 VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__nand4_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08324_ _01210_ _01223_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08255_ _01154_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08186_ _00547_ _00557_ _00556_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__a21bo_1
X_07206_ _02800_ _00109_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07137_ _05597_ _00040_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__nand2_1
X_07068_ _06380_ _06381_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__nor2_1
Xoutput261 net261 VGND VGND VPWR VPWR data_out[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput283 net283 VGND VGND VPWR VPWR data_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput272 net272 VGND VGND VPWR VPWR data_out[22] sky130_fd_sc_hd__clkbuf_4
X_09709_ _02584_ _02650_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__nor3_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10981_ _06416_ _00438_ net109 _02164_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__and4_1
X_12720_ _05951_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12651_ _05854_ _05855_ _05877_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__nor3_1
XFILLER_0_65_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11602_ _04291_ _04258_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12582_ _05799_ _05616_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__o21ai_1
X_11533_ _04637_ _04652_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11464_ _00479_ _03499_ _04576_ _04577_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10415_ _03385_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__xnor2_1
X_11395_ _02765_ _04500_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__a21bo_1
X_10346_ _03347_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _03272_ _03273_ _03256_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12016_ _04773_ _04787_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12849_ _02174_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08040_ _00939_ net82 net68 _00938_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09991_ _02956_ _02277_ _02960_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08942_ _01840_ _01841_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08873_ _00648_ _01196_ _01194_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07824_ _00724_ _00725_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__nor2_1
X_07755_ _00639_ _00640_ _00656_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06706_ net184 VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__clkbuf_4
X_07686_ _00339_ _00340_ _00587_ _00588_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__or4bb_4
X_09425_ _02338_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__and2b_1
X_06637_ _04292_ _02240_ _04325_ _04347_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__nand4_4
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ _01616_ _01623_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06568_ _03579_ _02657_ _03590_ _02668_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__a22o_1
X_06499_ _02789_ _02800_ _02811_ _02822_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__and4_4
XFILLER_0_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09287_ _02186_ _02187_ _01537_ _01539_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__o211ai_2
X_08307_ _00694_ _00696_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08238_ _00799_ _00801_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08169_ _01069_ _01070_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__or2_1
X_10200_ _02526_ _02528_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11180_ _03746_ _03766_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10131_ _03112_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10062_ _03037_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10964_ net81 net74 net75 net80 VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__a22o_1
X_12703_ _05878_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__nor2_1
X_10895_ _03945_ _03951_ _03953_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12634_ _05858_ _05859_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12565_ _01872_ _03210_ _04869_ _05245_ _05551_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__a41o_1
XFILLER_0_93_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11516_ _04152_ _04159_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12496_ _05642_ _05709_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11447_ _04557_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11378_ _03961_ _04482_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10329_ _03324_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xor2_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ _00030_ _00441_ _00442_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__nand3_2
XFILLER_0_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07471_ _00372_ _00373_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09210_ _01549_ _01550_ _01698_ _01696_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09141_ net50 net66 net5 _02470_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09072_ _01969_ _01970_ _01767_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08023_ _00456_ _00923_ _00924_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09974_ _02891_ _02942_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__xnor2_1
X_08925_ _01220_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__xnor2_1
X_08856_ _01753_ _01755_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07807_ _00708_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__inv_2
X_08787_ _01626_ _01627_ _01686_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07738_ _00268_ _00279_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__and2b_1
X_07669_ _00569_ _00570_ _00529_ _00127_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__o211a_1
X_09408_ _01657_ _02320_ _02321_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__and3_1
X_10680_ _03715_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09339_ _02237_ _02244_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__nand3_2
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12350_ _05547_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11301_ _03867_ _03868_ _03870_ _03871_ _03866_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12281_ _04762_ _05118_ _05117_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11232_ _00672_ _01835_ _04320_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11163_ _02185_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10114_ net170 net162 _01188_ net169 VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__a22o_1
X_11094_ _00543_ net48 VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__nand2_1
X_10045_ _03106_ net12 net223 net234 VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11996_ _01157_ _02464_ _05159_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10947_ _03986_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10878_ _03922_ _03934_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__xor2_4
XFILLER_0_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12617_ _05694_ _05840_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12548_ _05752_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__xnor2_1
XANTENNA_2 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12479_ _02215_ _03499_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _02229_ _06283_ _06284_ _02240_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ net211 net205 VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__and2_1
X_08710_ _04752_ _00516_ _01609_ _01610_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__nand4_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08641_ _00463_ _00964_ _01541_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08572_ _01470_ _01471_ _03579_ net82 VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__and4bb_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07523_ _06423_ _00420_ _00424_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__nor3_1
X_07454_ net2 VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07385_ _00264_ _00265_ _00286_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o21ba_1
X_09124_ _05882_ _06375_ _06368_ _00357_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09055_ _01934_ _01935_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08006_ _00452_ _00465_ _00907_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap293 _02579_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__buf_1
X_09957_ _02923_ _02924_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__nand2_2
X_08908_ _06254_ net91 net92 _04413_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__a22o_1
X_09888_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__inv_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _01737_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nor2_1
X_11850_ _04985_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__xor2_4
X_10801_ _03254_ _03303_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__a21o_1
X_11781_ _04923_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10732_ _03163_ _03770_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10663_ _03313_ _03129_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10594_ _04939_ _00549_ net56 net67 VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__and4_2
X_12402_ _05605_ _03967_ _04948_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12333_ _04781_ _05189_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12264_ _05053_ _05099_ _05454_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11215_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12195_ _05369_ _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11146_ _03671_ _03673_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nor2_1
X_11077_ net49 VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__buf_2
Xinput161 data_in[244] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xinput172 data_in[254] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
Xinput150 data_in[234] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
X_10028_ _02331_ _02333_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput183 data_in[33] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xinput194 data_in[43] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11979_ _02185_ _05141_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07170_ _00072_ _00073_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09811_ _02754_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__xnor2_2
X_09742_ net247 net239 net248 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06954_ _06265_ _06266_ _06140_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__a21oi_1
X_09673_ _01904_ _01907_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nand2_1
X_06885_ _06197_ _06198_ _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__a21oi_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ net100 net177 net178 net89 VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__a22o_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _00425_ _00946_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__and2_1
X_07506_ _06357_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__inv_2
X_08486_ _03864_ net240 net241 _02492_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07437_ _00337_ _00338_ _00193_ _00194_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07368_ _04238_ _06243_ _00270_ _02317_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__a22o_1
X_09107_ _05980_ _00830_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07299_ _04303_ _06283_ _00201_ _02229_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09038_ _06177_ net153 net154 net140 VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11000_ _04065_ _04066_ _04067_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11902_ _05056_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__xor2_4
XFILLER_0_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12882_ clknet_1_0__leaf_clk _00006_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dfxtp_1
X_11833_ _04978_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04893_ _04904_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _04365_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10715_ _06261_ net31 _03752_ _03753_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _03076_ _03077_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer5 _00600_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10577_ net37 net46 net38 net47 VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _05510_ _05507_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__or2b_1
X_12247_ _05435_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12178_ _05359_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__or2_1
X_11129_ _04136_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06670_ _04710_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08340_ _00716_ _00726_ _00724_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08271_ _01139_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07222_ _00123_ _00124_ _00106_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07153_ _00055_ _00056_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07084_ _06396_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07986_ _00885_ _00886_ _00393_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__a21bo_1
X_09725_ _01996_ _01999_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__nand2_2
X_06937_ _06249_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__xnor2_2
X_09656_ _02590_ _02593_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06868_ _06179_ _06180_ _06181_ _06176_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _01505_ _01506_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__nand3_4
X_09587_ _01234_ _01815_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__and2_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06799_ _05860_ _06104_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__and2_1
X_08538_ _01433_ _01437_ _01438_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08469_ _01364_ _01369_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10500_ _02940_ _02939_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__or2b_1
X_11480_ _04533_ _04535_ _04594_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10431_ _03437_ _03442_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10362_ _03366_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10293_ _06173_ _06304_ net206 net207 VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__and4_1
X_12101_ _04975_ _05023_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__a21o_1
X_12032_ _00672_ _03180_ _04800_ _04798_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12865_ _06103_ _02174_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__and3b_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _05970_ _05972_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11816_ _04942_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__xor2_2
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11747_ _04765_ _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__xor2_4
XFILLER_0_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11678_ _04805_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10629_ _03519_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07840_ net150 net142 net151 net141 VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ net94 _00672_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__nand2_1
X_09510_ _02431_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__and2_1
X_06722_ _03436_ _05279_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09441_ _02337_ _02356_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06653_ _04391_ _04402_ _04512_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__a21oi_1
X_09372_ net32 net48 _01632_ _01631_ _00530_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06584_ _03754_ _03765_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08323_ _01210_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08254_ _00620_ _01153_ _01152_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__a21oi_1
X_08185_ _01084_ _01085_ _01077_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__a21o_1
X_07205_ net23 VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__buf_2
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07136_ _06409_ _00039_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__xnor2_1
X_07067_ _06379_ _06378_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput262 net262 VGND VGND VPWR VPWR data_out[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput284 net284 VGND VGND VPWR VPWR data_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput273 net273 VGND VGND VPWR VPWR data_out[23] sky130_fd_sc_hd__clkbuf_4
X_09708_ _02648_ _02649_ _02000_ _02585_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__a211oi_2
X_07969_ _00388_ _00390_ _00389_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__a21bo_1
X_10980_ _00438_ _01520_ _02164_ _06416_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a22oi_2
X_09639_ _02542_ _02574_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12650_ _05854_ _05855_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11601_ _04243_ _04247_ _04726_ _04722_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__a31o_1
X_12581_ _05800_ _05801_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11532_ _04637_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11463_ _04573_ _04574_ _04575_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__nand3_1
X_10414_ _03422_ _03424_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11394_ _00872_ net57 net58 _00397_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__a22o_1
X_10345_ net254 net14 VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10276_ _03256_ _03272_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__and3_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _04788_ _04771_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__or2b_1
Xmax_cap3 _00149_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12848_ _06079_ _06084_ _06080_ net271 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__or4b_4
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12779_ _06014_ _06017_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _02957_ _02958_ _02959_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08941_ _01212_ _01214_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__or2_1
X_08872_ _01240_ _01241_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor2_1
X_07823_ _00205_ _00723_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07754_ _00259_ _00655_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__xor2_1
X_06705_ net183 _03348_ net184 _02712_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__a22o_1
X_07685_ _00585_ _00586_ _00143_ _00145_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__o211ai_1
X_09424_ _00109_ _00550_ _00544_ _00549_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a22o_1
X_06636_ _02229_ _04336_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_4
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09355_ _02261_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nor2_2
X_06567_ net77 VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06498_ _02789_ _02800_ _02811_ _02822_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a22oi_4
X_08306_ _00709_ _01206_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__xnor2_1
X_09286_ _01537_ _01539_ _02186_ _02187_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08237_ net303 _00632_ _00630_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08168_ _02811_ _01068_ _00545_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08099_ _00984_ _01000_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__xnor2_1
X_07119_ _06414_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10130_ _02431_ _02436_ _03111_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10061_ _02302_ _02366_ _03038_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10963_ net80 net81 net74 VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12702_ _05853_ _05880_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__and2b_1
X_10894_ _03949_ _03950_ _03946_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12633_ _03967_ _04948_ _05298_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a21oi_1
X_12564_ _05546_ _05556_ _05782_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11515_ _04156_ _04158_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12495_ _05705_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11446_ _06416_ _01520_ _04558_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21o_1
X_11377_ _03962_ _03969_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10328_ _02676_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _02601_ _02604_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07470_ _05980_ net246 _00370_ _00371_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _02038_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09071_ _01767_ _01969_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08022_ _03524_ _00438_ _00921_ _00922_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__nand4_2
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09973_ _02925_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08924_ _01822_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__nor2_1
X_08855_ _02328_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__and2_1
X_08786_ _01684_ _01685_ _01093_ net324 VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__a211o_1
X_07806_ net24 net25 _00239_ _00706_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__and4_1
X_07737_ _00269_ _00276_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07668_ _00529_ _00127_ net302 _00570_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09407_ _02318_ _02319_ _02309_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__a21o_1
X_06619_ _04128_ _02383_ _04139_ _02394_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a22o_1
X_07599_ _00072_ _00501_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__or2_1
X_09338_ _02242_ _02243_ _01605_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11300_ _03881_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__xnor2_1
X_09269_ net89 net100 _00453_ _00953_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12280_ _05178_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11231_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11162_ _03691_ _03692_ _04245_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10113_ _02427_ _02425_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__or2b_1
X_11093_ _04169_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10044_ net12 _01667_ _03019_ _03106_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11995_ _01157_ _05159_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10946_ _03987_ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10877_ _03924_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__xnor2_4
X_12616_ _05436_ _05692_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12547_ _05754_ _05764_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__xnor2_1
X_12478_ _05376_ _05372_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__and2b_1
XANTENNA_3 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11429_ _04538_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ net88 VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__clkbuf_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _00963_ _00952_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__or2b_1
X_08571_ _03579_ _00937_ _01470_ _01471_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07522_ _06423_ _00420_ _00424_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__o21a_1
X_07453_ _06373_ _00355_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09123_ _02481_ _02019_ _02020_ _02021_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__nand4_2
XFILLER_0_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07384_ _00264_ _00265_ _00286_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09054_ _01936_ _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08005_ _00031_ _00464_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap294 _01103_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09956_ _02920_ _02922_ _02903_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__a21o_1
X_08907_ _01231_ _01233_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__nand2_1
X_09887_ _02815_ _02153_ _02846_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__o211a_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _06243_ _06227_ _00270_ _00171_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__and4_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08769_ _01665_ _01668_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__nand3_1
X_10800_ _03305_ _03253_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__and2b_1
X_11780_ _00879_ _03967_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10731_ _03771_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__or2_1
X_12401_ _02765_ _03967_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10662_ _03086_ _03122_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__a21bo_2
X_10593_ _00549_ net56 net67 _04939_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12332_ _05523_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12263_ _05096_ _05098_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11214_ net29 _01217_ _01181_ net20 VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a22o_1
X_12194_ _05370_ _05377_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__xor2_1
X_11145_ _03739_ _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11076_ _00107_ _01629_ _03606_ _03605_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a31o_1
Xinput162 data_in[245] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
Xinput151 data_in[235] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xinput140 data_in[225] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_2
X_10027_ _02980_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__xnor2_4
Xinput173 data_in[255] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
Xinput184 data_in[34] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_4
Xinput195 data_in[44] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11978_ _04727_ _05140_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__or2_1
X_10929_ _00387_ net65 _03989_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09810_ _02761_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09741_ _02670_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__xor2_4
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06953_ _06140_ _06265_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09672_ _01927_ _01928_ _01929_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__nand3_1
XFILLER_0_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06884_ _04216_ _04589_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08623_ net180 VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_4
X_08554_ _01442_ _01454_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__xor2_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07505_ _00406_ _00407_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08485_ _02492_ _03864_ _00834_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07436_ _00193_ _00194_ _00337_ _00338_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_134_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07367_ net161 VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_4
X_09106_ _00834_ _02004_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09037_ _00775_ _01314_ _01313_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__a21o_1
X_07298_ net135 VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09939_ _05115_ _01562_ _02904_ _03337_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a22oi_1
X_11901_ _01667_ _01652_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12881_ clknet_1_0__leaf_clk _00005_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dfxtp_1
X_11832_ _04553_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__xnor2_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _04893_ _04904_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _04827_ _04828_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10714_ _06261_ _01784_ _03752_ _03753_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__a22oi_2
X_10645_ _03079_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10576_ _00530_ _01068_ _01051_ _00543_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer6 _00579_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_1
X_12315_ _05507_ _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12246_ _01584_ _01562_ _02239_ _02904_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__and4_1
X_12177_ _05355_ _05357_ _05358_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a21oi_1
X_11128_ _04207_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11059_ _04121_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08270_ _01169_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07221_ _00106_ _00123_ _00124_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07152_ _00053_ _00054_ _05158_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07083_ _06367_ _06395_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07985_ _00393_ _00885_ _00886_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__nand3b_1
X_09724_ _02192_ _02194_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__nand2_2
X_06936_ _02207_ _06142_ _04468_ _06145_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__a31o_1
X_09655_ _04128_ _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nand2_1
X_06867_ _06176_ _06179_ _06180_ _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__and4_1
X_08606_ _00920_ _00926_ _00925_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__a21bo_1
X_09586_ _01806_ _01814_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _05860_ _06104_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__nor2_1
X_08537_ _02580_ _01434_ _01435_ _01436_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__nand4_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ _01366_ _01368_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07419_ _00320_ _00321_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08399_ _01297_ _01298_ _01292_ _01294_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__a211o_1
X_10430_ _03440_ _03441_ _02817_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10361_ net8 net9 net4 net5 VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10292_ _06304_ _01365_ _01986_ _06173_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__a22oi_1
X_12100_ _04977_ _05022_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12031_ _05183_ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12864_ _06102_ _06100_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand2_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _05966_ _05968_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__or2_1
X_11815_ _04944_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__xor2_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11746_ _04842_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__xor2_4
XFILLER_0_56_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11677_ _04806_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__xnor2_1
X_10628_ _03658_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__xor2_4
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10559_ _02957_ _02959_ _02958_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12229_ _05416_ _04154_ _05068_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07770_ net91 VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__buf_2
X_06721_ _05180_ _05268_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__xor2_1
X_09440_ _02353_ _02354_ _02355_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06652_ _04391_ _04402_ _04512_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__and3_1
X_09371_ _02272_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__xnor2_1
X_06583_ _03732_ _02569_ _03743_ _02580_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08322_ _00710_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08253_ _00620_ _01152_ _01153_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__and3_1
X_07204_ _02800_ _03128_ _04972_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08184_ _01077_ _01084_ _01085_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07135_ _00037_ _00038_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07066_ _06378_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 net285 VGND VGND VPWR VPWR data_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput263 net263 VGND VGND VPWR VPWR data_out[14] sky130_fd_sc_hd__clkbuf_4
Xoutput274 net274 VGND VGND VPWR VPWR data_out[24] sky130_fd_sc_hd__clkbuf_4
X_07968_ _00386_ _00393_ _00394_ _00396_ _00400_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__a32o_1
X_09707_ _02000_ _02585_ _02648_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__o211a_1
X_06919_ _04490_ _06132_ _06231_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07899_ _00638_ _00799_ _00800_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__nor3_1
X_09638_ _02572_ _02573_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09569_ net22 VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__buf_2
X_12580_ _03859_ _05253_ _05569_ _05571_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__o2bb2ai_4
X_11600_ net260 _04720_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11531_ _04646_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11462_ _04573_ _04574_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11393_ _00397_ _00872_ _01444_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__and3_1
X_10413_ _02750_ _02784_ _03423_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__a21oi_2
X_10344_ _06375_ _00357_ net11 net13 VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10275_ _03269_ _03270_ _03262_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _04892_ _04969_ _04971_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap4 _01103_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_1
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ net271 _06087_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__or2b_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _06015_ _05950_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a21oi_1
X_11729_ _00810_ _02626_ _04409_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08940_ _01838_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__nor2_1
X_08871_ _00651_ _01198_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__nor2_1
X_07822_ _00205_ _00723_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07753_ _00278_ _00654_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06704_ net193 VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07684_ _00143_ _00145_ _00585_ _00586_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__a211o_1
X_09423_ net190 net23 _00550_ net34 VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06635_ _04303_ _02218_ _04314_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__and3_2
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09354_ _02259_ _02260_ _02200_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06566_ net69 VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08305_ _01204_ _01205_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06497_ net32 VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09285_ _02183_ _02184_ _02159_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08236_ _00637_ _01117_ _01118_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__nand3_2
X_08167_ net41 _01068_ _00545_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__and3_1
X_07118_ _06415_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__xor2_1
X_08098_ _00998_ _00999_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__nor2_1
X_07049_ _02448_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10060_ _01682_ _01684_ _02363_ _02364_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10962_ _03466_ _03474_ _03473_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_97_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12701_ _05796_ _05812_ _05810_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a21o_1
X_10893_ _03946_ _03949_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12632_ _03967_ _04948_ _05298_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__and3_2
XFILLER_0_136_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12563_ _05552_ _05554_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11514_ _04603_ _04632_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__xor2_4
XFILLER_0_81_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12494_ _05388_ _05457_ _05706_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11445_ _00438_ _02164_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11376_ _03962_ _03969_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10327_ _03325_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__xor2_4
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _02670_ _02685_ _02684_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a21o_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ _02504_ _02506_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09070_ _01967_ _01968_ _01768_ _01769_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08021_ _03524_ _00438_ _00921_ _00922_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09972_ _02939_ _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__xor2_2
XFILLER_0_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08923_ _01820_ _01821_ _06261_ net28 VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08854_ net173 VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__buf_4
X_08785_ _01093_ net300 _01684_ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_98_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07805_ _04446_ _00239_ _00706_ _02196_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a22o_1
X_07736_ _06331_ _00331_ _00335_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07667_ _00567_ _00568_ _00542_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09406_ _02309_ _02318_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__nand3_1
X_06618_ _04128_ _02383_ _04139_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__and3_1
X_07598_ _00093_ _00500_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09337_ _01605_ _02242_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__nand3_2
XFILLER_0_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06549_ net174 VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09268_ _02163_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__xor2_2
XFILLER_0_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08219_ _00591_ _00593_ _01119_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ _02059_ _02097_ _02098_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__nand3_1
X_11230_ net98 net99 net92 net93 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11161_ _03691_ _03692_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10112_ _02424_ _02419_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__or2b_1
X_11092_ net46 net38 net47 net39 VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__and4_1
X_10043_ net234 VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11994_ _00617_ _02464_ _03709_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__and3_1
X_10945_ _03997_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__xor2_2
X_10876_ _03925_ _03932_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12615_ _05690_ _05697_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12546_ _05762_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12477_ _05370_ _05377_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nand2_1
X_11428_ _00421_ net82 _01488_ net75 VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__and4_2
XANTENNA_4 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11359_ _00357_ _02019_ _04460_ _04461_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__nand4_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08570_ net70 net71 net80 net81 VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07521_ _00422_ _00423_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ net6 net7 net255 net2 VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ _00284_ _00285_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09122_ net252 _02019_ _02020_ _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09053_ _01951_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08004_ _00903_ _00904_ _00806_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap295 _00792_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09955_ _02903_ _02920_ _02922_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__nand3_2
X_08906_ _01252_ _01253_ _01261_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__o31a_1
X_09886_ _02843_ _02845_ _02829_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__o21ai_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08837_ _06227_ _00270_ _00171_ _06243_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__a22oi_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _03106_ net212 net223 _02789_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08699_ _01598_ _01597_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__or2b_1
X_07719_ _00273_ _00275_ _00619_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o21a_1
X_10730_ _06264_ _00250_ _01217_ _02498_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10661_ _03089_ _03121_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12400_ _04949_ _05308_ _04951_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10592_ _00549_ net45 _03015_ _03014_ _01666_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12331_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12262_ _05430_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11213_ _03777_ _03792_ _03791_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12193_ _05372_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11144_ _04224_ _04226_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__xor2_2
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11075_ _04145_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput152 data_in[236] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
Xinput141 data_in[226] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
Xinput130 data_in[216] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
Xinput163 data_in[246] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
X_10026_ _02999_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__or2b_2
Xinput174 data_in[25] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
Xinput196 data_in[45] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
Xinput185 data_in[35] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11977_ _04727_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__nand2_1
X_10928_ net63 net55 net64 net57 VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__nand4_2
XFILLER_0_39_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10859_ _03741_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12529_ _02174_ _05744_ _05745_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09740_ _02684_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__or2b_2
X_06952_ _04435_ _06142_ _06264_ _02207_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__a22o_1
.ends

