magic
tech sky130A
magscale 1 2
timestamp 1695331800
<< obsli1 >>
rect 1104 2159 75808 76721
<< obsm1 >>
rect 1104 1912 75886 77648
<< metal2 >>
rect 3238 78308 3294 79108
rect 3514 78308 3570 79108
rect 3790 78308 3846 79108
rect 4066 78308 4122 79108
rect 4342 78308 4398 79108
rect 4618 78308 4674 79108
rect 4894 78308 4950 79108
rect 5170 78308 5226 79108
rect 5446 78308 5502 79108
rect 5722 78308 5778 79108
rect 5998 78308 6054 79108
rect 6274 78308 6330 79108
rect 6550 78308 6606 79108
rect 6826 78308 6882 79108
rect 7102 78308 7158 79108
rect 7378 78308 7434 79108
rect 7654 78308 7710 79108
rect 7930 78308 7986 79108
rect 8206 78308 8262 79108
rect 8482 78308 8538 79108
rect 8758 78308 8814 79108
rect 9034 78308 9090 79108
rect 9310 78308 9366 79108
rect 9586 78308 9642 79108
rect 9862 78308 9918 79108
rect 10138 78308 10194 79108
rect 10414 78308 10470 79108
rect 10690 78308 10746 79108
rect 10966 78308 11022 79108
rect 11242 78308 11298 79108
rect 11518 78308 11574 79108
rect 11794 78308 11850 79108
rect 12070 78308 12126 79108
rect 12346 78308 12402 79108
rect 12622 78308 12678 79108
rect 12898 78308 12954 79108
rect 13174 78308 13230 79108
rect 13450 78308 13506 79108
rect 13726 78308 13782 79108
rect 14002 78308 14058 79108
rect 14278 78308 14334 79108
rect 14554 78308 14610 79108
rect 14830 78308 14886 79108
rect 15106 78308 15162 79108
rect 15382 78308 15438 79108
rect 15658 78308 15714 79108
rect 15934 78308 15990 79108
rect 16210 78308 16266 79108
rect 16486 78308 16542 79108
rect 16762 78308 16818 79108
rect 17038 78308 17094 79108
rect 17314 78308 17370 79108
rect 17590 78308 17646 79108
rect 17866 78308 17922 79108
rect 18142 78308 18198 79108
rect 18418 78308 18474 79108
rect 18694 78308 18750 79108
rect 18970 78308 19026 79108
rect 19246 78308 19302 79108
rect 19522 78308 19578 79108
rect 19798 78308 19854 79108
rect 20074 78308 20130 79108
rect 20350 78308 20406 79108
rect 20626 78308 20682 79108
rect 20902 78308 20958 79108
rect 21178 78308 21234 79108
rect 21454 78308 21510 79108
rect 21730 78308 21786 79108
rect 22006 78308 22062 79108
rect 22282 78308 22338 79108
rect 22558 78308 22614 79108
rect 22834 78308 22890 79108
rect 23110 78308 23166 79108
rect 23386 78308 23442 79108
rect 23662 78308 23718 79108
rect 23938 78308 23994 79108
rect 24214 78308 24270 79108
rect 24490 78308 24546 79108
rect 24766 78308 24822 79108
rect 25042 78308 25098 79108
rect 25318 78308 25374 79108
rect 25594 78308 25650 79108
rect 25870 78308 25926 79108
rect 26146 78308 26202 79108
rect 26422 78308 26478 79108
rect 26698 78308 26754 79108
rect 26974 78308 27030 79108
rect 27250 78308 27306 79108
rect 27526 78308 27582 79108
rect 27802 78308 27858 79108
rect 28078 78308 28134 79108
rect 28354 78308 28410 79108
rect 28630 78308 28686 79108
rect 28906 78308 28962 79108
rect 29182 78308 29238 79108
rect 29458 78308 29514 79108
rect 29734 78308 29790 79108
rect 30010 78308 30066 79108
rect 30286 78308 30342 79108
rect 30562 78308 30618 79108
rect 30838 78308 30894 79108
rect 31114 78308 31170 79108
rect 31390 78308 31446 79108
rect 31666 78308 31722 79108
rect 31942 78308 31998 79108
rect 32218 78308 32274 79108
rect 32494 78308 32550 79108
rect 32770 78308 32826 79108
rect 33046 78308 33102 79108
rect 33322 78308 33378 79108
rect 33598 78308 33654 79108
rect 33874 78308 33930 79108
rect 34150 78308 34206 79108
rect 34426 78308 34482 79108
rect 34702 78308 34758 79108
rect 34978 78308 35034 79108
rect 35254 78308 35310 79108
rect 35530 78308 35586 79108
rect 35806 78308 35862 79108
rect 36082 78308 36138 79108
rect 36358 78308 36414 79108
rect 36634 78308 36690 79108
rect 36910 78308 36966 79108
rect 37186 78308 37242 79108
rect 37462 78308 37518 79108
rect 37738 78308 37794 79108
rect 38014 78308 38070 79108
rect 38290 78308 38346 79108
rect 38566 78308 38622 79108
rect 38842 78308 38898 79108
rect 39118 78308 39174 79108
rect 39394 78308 39450 79108
rect 39670 78308 39726 79108
rect 39946 78308 40002 79108
rect 40222 78308 40278 79108
rect 40498 78308 40554 79108
rect 40774 78308 40830 79108
rect 41050 78308 41106 79108
rect 41326 78308 41382 79108
rect 41602 78308 41658 79108
rect 41878 78308 41934 79108
rect 42154 78308 42210 79108
rect 42430 78308 42486 79108
rect 42706 78308 42762 79108
rect 42982 78308 43038 79108
rect 43258 78308 43314 79108
rect 43534 78308 43590 79108
rect 43810 78308 43866 79108
rect 44086 78308 44142 79108
rect 44362 78308 44418 79108
rect 44638 78308 44694 79108
rect 44914 78308 44970 79108
rect 45190 78308 45246 79108
rect 45466 78308 45522 79108
rect 45742 78308 45798 79108
rect 46018 78308 46074 79108
rect 46294 78308 46350 79108
rect 46570 78308 46626 79108
rect 46846 78308 46902 79108
rect 47122 78308 47178 79108
rect 47398 78308 47454 79108
rect 47674 78308 47730 79108
rect 47950 78308 48006 79108
rect 48226 78308 48282 79108
rect 48502 78308 48558 79108
rect 48778 78308 48834 79108
rect 49054 78308 49110 79108
rect 49330 78308 49386 79108
rect 49606 78308 49662 79108
rect 49882 78308 49938 79108
rect 50158 78308 50214 79108
rect 50434 78308 50490 79108
rect 50710 78308 50766 79108
rect 50986 78308 51042 79108
rect 51262 78308 51318 79108
rect 51538 78308 51594 79108
rect 51814 78308 51870 79108
rect 52090 78308 52146 79108
rect 52366 78308 52422 79108
rect 52642 78308 52698 79108
rect 52918 78308 52974 79108
rect 53194 78308 53250 79108
rect 53470 78308 53526 79108
rect 53746 78308 53802 79108
rect 54022 78308 54078 79108
rect 54298 78308 54354 79108
rect 54574 78308 54630 79108
rect 54850 78308 54906 79108
rect 55126 78308 55182 79108
rect 55402 78308 55458 79108
rect 55678 78308 55734 79108
rect 55954 78308 56010 79108
rect 56230 78308 56286 79108
rect 56506 78308 56562 79108
rect 56782 78308 56838 79108
rect 57058 78308 57114 79108
rect 57334 78308 57390 79108
rect 57610 78308 57666 79108
rect 57886 78308 57942 79108
rect 58162 78308 58218 79108
rect 58438 78308 58494 79108
rect 58714 78308 58770 79108
rect 58990 78308 59046 79108
rect 59266 78308 59322 79108
rect 59542 78308 59598 79108
rect 59818 78308 59874 79108
rect 60094 78308 60150 79108
rect 60370 78308 60426 79108
rect 60646 78308 60702 79108
rect 60922 78308 60978 79108
rect 61198 78308 61254 79108
rect 61474 78308 61530 79108
rect 61750 78308 61806 79108
rect 62026 78308 62082 79108
rect 62302 78308 62358 79108
rect 62578 78308 62634 79108
rect 62854 78308 62910 79108
rect 63130 78308 63186 79108
rect 63406 78308 63462 79108
rect 63682 78308 63738 79108
rect 63958 78308 64014 79108
rect 64234 78308 64290 79108
rect 64510 78308 64566 79108
rect 64786 78308 64842 79108
rect 65062 78308 65118 79108
rect 65338 78308 65394 79108
rect 65614 78308 65670 79108
rect 65890 78308 65946 79108
rect 66166 78308 66222 79108
rect 66442 78308 66498 79108
rect 66718 78308 66774 79108
rect 66994 78308 67050 79108
rect 67270 78308 67326 79108
rect 67546 78308 67602 79108
rect 67822 78308 67878 79108
rect 68098 78308 68154 79108
rect 68374 78308 68430 79108
rect 68650 78308 68706 79108
rect 68926 78308 68982 79108
rect 69202 78308 69258 79108
rect 69478 78308 69534 79108
rect 69754 78308 69810 79108
rect 70030 78308 70086 79108
rect 70306 78308 70362 79108
rect 70582 78308 70638 79108
rect 70858 78308 70914 79108
rect 71134 78308 71190 79108
rect 71410 78308 71466 79108
rect 71686 78308 71742 79108
rect 71962 78308 72018 79108
rect 72238 78308 72294 79108
rect 72514 78308 72570 79108
rect 72790 78308 72846 79108
rect 73066 78308 73122 79108
rect 73342 78308 73398 79108
rect 73618 78308 73674 79108
rect 2410 0 2466 800
rect 5078 0 5134 800
rect 7746 0 7802 800
rect 10414 0 10470 800
rect 13082 0 13138 800
rect 15750 0 15806 800
rect 18418 0 18474 800
rect 21086 0 21142 800
rect 23754 0 23810 800
rect 26422 0 26478 800
rect 29090 0 29146 800
rect 31758 0 31814 800
rect 34426 0 34482 800
rect 37094 0 37150 800
rect 39762 0 39818 800
rect 42430 0 42486 800
rect 45098 0 45154 800
rect 47766 0 47822 800
rect 50434 0 50490 800
rect 53102 0 53158 800
rect 55770 0 55826 800
rect 58438 0 58494 800
rect 61106 0 61162 800
rect 63774 0 63830 800
rect 66442 0 66498 800
rect 69110 0 69166 800
rect 71778 0 71834 800
rect 74446 0 74502 800
<< obsm2 >>
rect 1398 78252 3182 78418
rect 3350 78252 3458 78418
rect 3626 78252 3734 78418
rect 3902 78252 4010 78418
rect 4178 78252 4286 78418
rect 4454 78252 4562 78418
rect 4730 78252 4838 78418
rect 5006 78252 5114 78418
rect 5282 78252 5390 78418
rect 5558 78252 5666 78418
rect 5834 78252 5942 78418
rect 6110 78252 6218 78418
rect 6386 78252 6494 78418
rect 6662 78252 6770 78418
rect 6938 78252 7046 78418
rect 7214 78252 7322 78418
rect 7490 78252 7598 78418
rect 7766 78252 7874 78418
rect 8042 78252 8150 78418
rect 8318 78252 8426 78418
rect 8594 78252 8702 78418
rect 8870 78252 8978 78418
rect 9146 78252 9254 78418
rect 9422 78252 9530 78418
rect 9698 78252 9806 78418
rect 9974 78252 10082 78418
rect 10250 78252 10358 78418
rect 10526 78252 10634 78418
rect 10802 78252 10910 78418
rect 11078 78252 11186 78418
rect 11354 78252 11462 78418
rect 11630 78252 11738 78418
rect 11906 78252 12014 78418
rect 12182 78252 12290 78418
rect 12458 78252 12566 78418
rect 12734 78252 12842 78418
rect 13010 78252 13118 78418
rect 13286 78252 13394 78418
rect 13562 78252 13670 78418
rect 13838 78252 13946 78418
rect 14114 78252 14222 78418
rect 14390 78252 14498 78418
rect 14666 78252 14774 78418
rect 14942 78252 15050 78418
rect 15218 78252 15326 78418
rect 15494 78252 15602 78418
rect 15770 78252 15878 78418
rect 16046 78252 16154 78418
rect 16322 78252 16430 78418
rect 16598 78252 16706 78418
rect 16874 78252 16982 78418
rect 17150 78252 17258 78418
rect 17426 78252 17534 78418
rect 17702 78252 17810 78418
rect 17978 78252 18086 78418
rect 18254 78252 18362 78418
rect 18530 78252 18638 78418
rect 18806 78252 18914 78418
rect 19082 78252 19190 78418
rect 19358 78252 19466 78418
rect 19634 78252 19742 78418
rect 19910 78252 20018 78418
rect 20186 78252 20294 78418
rect 20462 78252 20570 78418
rect 20738 78252 20846 78418
rect 21014 78252 21122 78418
rect 21290 78252 21398 78418
rect 21566 78252 21674 78418
rect 21842 78252 21950 78418
rect 22118 78252 22226 78418
rect 22394 78252 22502 78418
rect 22670 78252 22778 78418
rect 22946 78252 23054 78418
rect 23222 78252 23330 78418
rect 23498 78252 23606 78418
rect 23774 78252 23882 78418
rect 24050 78252 24158 78418
rect 24326 78252 24434 78418
rect 24602 78252 24710 78418
rect 24878 78252 24986 78418
rect 25154 78252 25262 78418
rect 25430 78252 25538 78418
rect 25706 78252 25814 78418
rect 25982 78252 26090 78418
rect 26258 78252 26366 78418
rect 26534 78252 26642 78418
rect 26810 78252 26918 78418
rect 27086 78252 27194 78418
rect 27362 78252 27470 78418
rect 27638 78252 27746 78418
rect 27914 78252 28022 78418
rect 28190 78252 28298 78418
rect 28466 78252 28574 78418
rect 28742 78252 28850 78418
rect 29018 78252 29126 78418
rect 29294 78252 29402 78418
rect 29570 78252 29678 78418
rect 29846 78252 29954 78418
rect 30122 78252 30230 78418
rect 30398 78252 30506 78418
rect 30674 78252 30782 78418
rect 30950 78252 31058 78418
rect 31226 78252 31334 78418
rect 31502 78252 31610 78418
rect 31778 78252 31886 78418
rect 32054 78252 32162 78418
rect 32330 78252 32438 78418
rect 32606 78252 32714 78418
rect 32882 78252 32990 78418
rect 33158 78252 33266 78418
rect 33434 78252 33542 78418
rect 33710 78252 33818 78418
rect 33986 78252 34094 78418
rect 34262 78252 34370 78418
rect 34538 78252 34646 78418
rect 34814 78252 34922 78418
rect 35090 78252 35198 78418
rect 35366 78252 35474 78418
rect 35642 78252 35750 78418
rect 35918 78252 36026 78418
rect 36194 78252 36302 78418
rect 36470 78252 36578 78418
rect 36746 78252 36854 78418
rect 37022 78252 37130 78418
rect 37298 78252 37406 78418
rect 37574 78252 37682 78418
rect 37850 78252 37958 78418
rect 38126 78252 38234 78418
rect 38402 78252 38510 78418
rect 38678 78252 38786 78418
rect 38954 78252 39062 78418
rect 39230 78252 39338 78418
rect 39506 78252 39614 78418
rect 39782 78252 39890 78418
rect 40058 78252 40166 78418
rect 40334 78252 40442 78418
rect 40610 78252 40718 78418
rect 40886 78252 40994 78418
rect 41162 78252 41270 78418
rect 41438 78252 41546 78418
rect 41714 78252 41822 78418
rect 41990 78252 42098 78418
rect 42266 78252 42374 78418
rect 42542 78252 42650 78418
rect 42818 78252 42926 78418
rect 43094 78252 43202 78418
rect 43370 78252 43478 78418
rect 43646 78252 43754 78418
rect 43922 78252 44030 78418
rect 44198 78252 44306 78418
rect 44474 78252 44582 78418
rect 44750 78252 44858 78418
rect 45026 78252 45134 78418
rect 45302 78252 45410 78418
rect 45578 78252 45686 78418
rect 45854 78252 45962 78418
rect 46130 78252 46238 78418
rect 46406 78252 46514 78418
rect 46682 78252 46790 78418
rect 46958 78252 47066 78418
rect 47234 78252 47342 78418
rect 47510 78252 47618 78418
rect 47786 78252 47894 78418
rect 48062 78252 48170 78418
rect 48338 78252 48446 78418
rect 48614 78252 48722 78418
rect 48890 78252 48998 78418
rect 49166 78252 49274 78418
rect 49442 78252 49550 78418
rect 49718 78252 49826 78418
rect 49994 78252 50102 78418
rect 50270 78252 50378 78418
rect 50546 78252 50654 78418
rect 50822 78252 50930 78418
rect 51098 78252 51206 78418
rect 51374 78252 51482 78418
rect 51650 78252 51758 78418
rect 51926 78252 52034 78418
rect 52202 78252 52310 78418
rect 52478 78252 52586 78418
rect 52754 78252 52862 78418
rect 53030 78252 53138 78418
rect 53306 78252 53414 78418
rect 53582 78252 53690 78418
rect 53858 78252 53966 78418
rect 54134 78252 54242 78418
rect 54410 78252 54518 78418
rect 54686 78252 54794 78418
rect 54962 78252 55070 78418
rect 55238 78252 55346 78418
rect 55514 78252 55622 78418
rect 55790 78252 55898 78418
rect 56066 78252 56174 78418
rect 56342 78252 56450 78418
rect 56618 78252 56726 78418
rect 56894 78252 57002 78418
rect 57170 78252 57278 78418
rect 57446 78252 57554 78418
rect 57722 78252 57830 78418
rect 57998 78252 58106 78418
rect 58274 78252 58382 78418
rect 58550 78252 58658 78418
rect 58826 78252 58934 78418
rect 59102 78252 59210 78418
rect 59378 78252 59486 78418
rect 59654 78252 59762 78418
rect 59930 78252 60038 78418
rect 60206 78252 60314 78418
rect 60482 78252 60590 78418
rect 60758 78252 60866 78418
rect 61034 78252 61142 78418
rect 61310 78252 61418 78418
rect 61586 78252 61694 78418
rect 61862 78252 61970 78418
rect 62138 78252 62246 78418
rect 62414 78252 62522 78418
rect 62690 78252 62798 78418
rect 62966 78252 63074 78418
rect 63242 78252 63350 78418
rect 63518 78252 63626 78418
rect 63794 78252 63902 78418
rect 64070 78252 64178 78418
rect 64346 78252 64454 78418
rect 64622 78252 64730 78418
rect 64898 78252 65006 78418
rect 65174 78252 65282 78418
rect 65450 78252 65558 78418
rect 65726 78252 65834 78418
rect 66002 78252 66110 78418
rect 66278 78252 66386 78418
rect 66554 78252 66662 78418
rect 66830 78252 66938 78418
rect 67106 78252 67214 78418
rect 67382 78252 67490 78418
rect 67658 78252 67766 78418
rect 67934 78252 68042 78418
rect 68210 78252 68318 78418
rect 68486 78252 68594 78418
rect 68762 78252 68870 78418
rect 69038 78252 69146 78418
rect 69314 78252 69422 78418
rect 69590 78252 69698 78418
rect 69866 78252 69974 78418
rect 70142 78252 70250 78418
rect 70418 78252 70526 78418
rect 70694 78252 70802 78418
rect 70970 78252 71078 78418
rect 71246 78252 71354 78418
rect 71522 78252 71630 78418
rect 71798 78252 71906 78418
rect 72074 78252 72182 78418
rect 72350 78252 72458 78418
rect 72626 78252 72734 78418
rect 72902 78252 73010 78418
rect 73178 78252 73286 78418
rect 73454 78252 73562 78418
rect 73730 78252 75880 78418
rect 1398 856 75880 78252
rect 1398 734 2354 856
rect 2522 734 5022 856
rect 5190 734 7690 856
rect 7858 734 10358 856
rect 10526 734 13026 856
rect 13194 734 15694 856
rect 15862 734 18362 856
rect 18530 734 21030 856
rect 21198 734 23698 856
rect 23866 734 26366 856
rect 26534 734 29034 856
rect 29202 734 31702 856
rect 31870 734 34370 856
rect 34538 734 37038 856
rect 37206 734 39706 856
rect 39874 734 42374 856
rect 42542 734 45042 856
rect 45210 734 47710 856
rect 47878 734 50378 856
rect 50546 734 53046 856
rect 53214 734 55714 856
rect 55882 734 58382 856
rect 58550 734 61050 856
rect 61218 734 63718 856
rect 63886 734 66386 856
rect 66554 734 69054 856
rect 69222 734 71722 856
rect 71890 734 74390 856
rect 74558 734 75880 856
<< metal3 >>
rect 0 59032 800 59152
rect 0 19592 800 19712
<< obsm3 >>
rect 798 59232 75703 77621
rect 880 58952 75703 59232
rect 798 19792 75703 58952
rect 880 19512 75703 19792
rect 798 2143 75703 19512
<< metal4 >>
rect 2344 2128 2664 76752
rect 3004 2128 3324 76752
rect 33064 2128 33384 76752
rect 33724 2128 34044 76752
rect 63784 2128 64104 76752
rect 64444 2128 64764 76752
<< obsm4 >>
rect 6499 76832 74093 77485
rect 6499 13499 32984 76832
rect 33464 13499 33644 76832
rect 34124 13499 63704 76832
rect 64184 13499 64364 76832
rect 64844 13499 74093 76832
<< metal5 >>
rect 1056 65348 75856 65668
rect 1056 64688 75856 65008
rect 1056 34712 75856 35032
rect 1056 34052 75856 34372
rect 1056 4076 75856 4396
rect 1056 3416 75856 3736
<< obsm5 >>
rect 17780 74980 40548 75980
<< labels >>
rlabel metal4 s 3004 2128 3324 76752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 33724 2128 34044 76752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 64444 2128 64764 76752 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4076 75856 4396 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 34712 75856 35032 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 65348 75856 65668 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2344 2128 2664 76752 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 33064 2128 33384 76752 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 63784 2128 64104 76752 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3416 75856 3736 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 34052 75856 34372 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 64688 75856 65008 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 19592 800 19712 6 clk
port 3 nsew signal input
rlabel metal2 s 3238 78308 3294 79108 6 data_in[0]
port 4 nsew signal input
rlabel metal2 s 30838 78308 30894 79108 6 data_in[100]
port 5 nsew signal input
rlabel metal2 s 31114 78308 31170 79108 6 data_in[101]
port 6 nsew signal input
rlabel metal2 s 31390 78308 31446 79108 6 data_in[102]
port 7 nsew signal input
rlabel metal2 s 31666 78308 31722 79108 6 data_in[103]
port 8 nsew signal input
rlabel metal2 s 31942 78308 31998 79108 6 data_in[104]
port 9 nsew signal input
rlabel metal2 s 32218 78308 32274 79108 6 data_in[105]
port 10 nsew signal input
rlabel metal2 s 32494 78308 32550 79108 6 data_in[106]
port 11 nsew signal input
rlabel metal2 s 32770 78308 32826 79108 6 data_in[107]
port 12 nsew signal input
rlabel metal2 s 33046 78308 33102 79108 6 data_in[108]
port 13 nsew signal input
rlabel metal2 s 33322 78308 33378 79108 6 data_in[109]
port 14 nsew signal input
rlabel metal2 s 5998 78308 6054 79108 6 data_in[10]
port 15 nsew signal input
rlabel metal2 s 33598 78308 33654 79108 6 data_in[110]
port 16 nsew signal input
rlabel metal2 s 33874 78308 33930 79108 6 data_in[111]
port 17 nsew signal input
rlabel metal2 s 34150 78308 34206 79108 6 data_in[112]
port 18 nsew signal input
rlabel metal2 s 34426 78308 34482 79108 6 data_in[113]
port 19 nsew signal input
rlabel metal2 s 34702 78308 34758 79108 6 data_in[114]
port 20 nsew signal input
rlabel metal2 s 34978 78308 35034 79108 6 data_in[115]
port 21 nsew signal input
rlabel metal2 s 35254 78308 35310 79108 6 data_in[116]
port 22 nsew signal input
rlabel metal2 s 35530 78308 35586 79108 6 data_in[117]
port 23 nsew signal input
rlabel metal2 s 35806 78308 35862 79108 6 data_in[118]
port 24 nsew signal input
rlabel metal2 s 36082 78308 36138 79108 6 data_in[119]
port 25 nsew signal input
rlabel metal2 s 6274 78308 6330 79108 6 data_in[11]
port 26 nsew signal input
rlabel metal2 s 36358 78308 36414 79108 6 data_in[120]
port 27 nsew signal input
rlabel metal2 s 36634 78308 36690 79108 6 data_in[121]
port 28 nsew signal input
rlabel metal2 s 36910 78308 36966 79108 6 data_in[122]
port 29 nsew signal input
rlabel metal2 s 37186 78308 37242 79108 6 data_in[123]
port 30 nsew signal input
rlabel metal2 s 37462 78308 37518 79108 6 data_in[124]
port 31 nsew signal input
rlabel metal2 s 37738 78308 37794 79108 6 data_in[125]
port 32 nsew signal input
rlabel metal2 s 38014 78308 38070 79108 6 data_in[126]
port 33 nsew signal input
rlabel metal2 s 38290 78308 38346 79108 6 data_in[127]
port 34 nsew signal input
rlabel metal2 s 38566 78308 38622 79108 6 data_in[128]
port 35 nsew signal input
rlabel metal2 s 38842 78308 38898 79108 6 data_in[129]
port 36 nsew signal input
rlabel metal2 s 6550 78308 6606 79108 6 data_in[12]
port 37 nsew signal input
rlabel metal2 s 39118 78308 39174 79108 6 data_in[130]
port 38 nsew signal input
rlabel metal2 s 39394 78308 39450 79108 6 data_in[131]
port 39 nsew signal input
rlabel metal2 s 39670 78308 39726 79108 6 data_in[132]
port 40 nsew signal input
rlabel metal2 s 39946 78308 40002 79108 6 data_in[133]
port 41 nsew signal input
rlabel metal2 s 40222 78308 40278 79108 6 data_in[134]
port 42 nsew signal input
rlabel metal2 s 40498 78308 40554 79108 6 data_in[135]
port 43 nsew signal input
rlabel metal2 s 40774 78308 40830 79108 6 data_in[136]
port 44 nsew signal input
rlabel metal2 s 41050 78308 41106 79108 6 data_in[137]
port 45 nsew signal input
rlabel metal2 s 41326 78308 41382 79108 6 data_in[138]
port 46 nsew signal input
rlabel metal2 s 41602 78308 41658 79108 6 data_in[139]
port 47 nsew signal input
rlabel metal2 s 6826 78308 6882 79108 6 data_in[13]
port 48 nsew signal input
rlabel metal2 s 41878 78308 41934 79108 6 data_in[140]
port 49 nsew signal input
rlabel metal2 s 42154 78308 42210 79108 6 data_in[141]
port 50 nsew signal input
rlabel metal2 s 42430 78308 42486 79108 6 data_in[142]
port 51 nsew signal input
rlabel metal2 s 42706 78308 42762 79108 6 data_in[143]
port 52 nsew signal input
rlabel metal2 s 42982 78308 43038 79108 6 data_in[144]
port 53 nsew signal input
rlabel metal2 s 43258 78308 43314 79108 6 data_in[145]
port 54 nsew signal input
rlabel metal2 s 43534 78308 43590 79108 6 data_in[146]
port 55 nsew signal input
rlabel metal2 s 43810 78308 43866 79108 6 data_in[147]
port 56 nsew signal input
rlabel metal2 s 44086 78308 44142 79108 6 data_in[148]
port 57 nsew signal input
rlabel metal2 s 44362 78308 44418 79108 6 data_in[149]
port 58 nsew signal input
rlabel metal2 s 7102 78308 7158 79108 6 data_in[14]
port 59 nsew signal input
rlabel metal2 s 44638 78308 44694 79108 6 data_in[150]
port 60 nsew signal input
rlabel metal2 s 44914 78308 44970 79108 6 data_in[151]
port 61 nsew signal input
rlabel metal2 s 45190 78308 45246 79108 6 data_in[152]
port 62 nsew signal input
rlabel metal2 s 45466 78308 45522 79108 6 data_in[153]
port 63 nsew signal input
rlabel metal2 s 45742 78308 45798 79108 6 data_in[154]
port 64 nsew signal input
rlabel metal2 s 46018 78308 46074 79108 6 data_in[155]
port 65 nsew signal input
rlabel metal2 s 46294 78308 46350 79108 6 data_in[156]
port 66 nsew signal input
rlabel metal2 s 46570 78308 46626 79108 6 data_in[157]
port 67 nsew signal input
rlabel metal2 s 46846 78308 46902 79108 6 data_in[158]
port 68 nsew signal input
rlabel metal2 s 47122 78308 47178 79108 6 data_in[159]
port 69 nsew signal input
rlabel metal2 s 7378 78308 7434 79108 6 data_in[15]
port 70 nsew signal input
rlabel metal2 s 47398 78308 47454 79108 6 data_in[160]
port 71 nsew signal input
rlabel metal2 s 47674 78308 47730 79108 6 data_in[161]
port 72 nsew signal input
rlabel metal2 s 47950 78308 48006 79108 6 data_in[162]
port 73 nsew signal input
rlabel metal2 s 48226 78308 48282 79108 6 data_in[163]
port 74 nsew signal input
rlabel metal2 s 48502 78308 48558 79108 6 data_in[164]
port 75 nsew signal input
rlabel metal2 s 48778 78308 48834 79108 6 data_in[165]
port 76 nsew signal input
rlabel metal2 s 49054 78308 49110 79108 6 data_in[166]
port 77 nsew signal input
rlabel metal2 s 49330 78308 49386 79108 6 data_in[167]
port 78 nsew signal input
rlabel metal2 s 49606 78308 49662 79108 6 data_in[168]
port 79 nsew signal input
rlabel metal2 s 49882 78308 49938 79108 6 data_in[169]
port 80 nsew signal input
rlabel metal2 s 7654 78308 7710 79108 6 data_in[16]
port 81 nsew signal input
rlabel metal2 s 50158 78308 50214 79108 6 data_in[170]
port 82 nsew signal input
rlabel metal2 s 50434 78308 50490 79108 6 data_in[171]
port 83 nsew signal input
rlabel metal2 s 50710 78308 50766 79108 6 data_in[172]
port 84 nsew signal input
rlabel metal2 s 50986 78308 51042 79108 6 data_in[173]
port 85 nsew signal input
rlabel metal2 s 51262 78308 51318 79108 6 data_in[174]
port 86 nsew signal input
rlabel metal2 s 51538 78308 51594 79108 6 data_in[175]
port 87 nsew signal input
rlabel metal2 s 51814 78308 51870 79108 6 data_in[176]
port 88 nsew signal input
rlabel metal2 s 52090 78308 52146 79108 6 data_in[177]
port 89 nsew signal input
rlabel metal2 s 52366 78308 52422 79108 6 data_in[178]
port 90 nsew signal input
rlabel metal2 s 52642 78308 52698 79108 6 data_in[179]
port 91 nsew signal input
rlabel metal2 s 7930 78308 7986 79108 6 data_in[17]
port 92 nsew signal input
rlabel metal2 s 52918 78308 52974 79108 6 data_in[180]
port 93 nsew signal input
rlabel metal2 s 53194 78308 53250 79108 6 data_in[181]
port 94 nsew signal input
rlabel metal2 s 53470 78308 53526 79108 6 data_in[182]
port 95 nsew signal input
rlabel metal2 s 53746 78308 53802 79108 6 data_in[183]
port 96 nsew signal input
rlabel metal2 s 54022 78308 54078 79108 6 data_in[184]
port 97 nsew signal input
rlabel metal2 s 54298 78308 54354 79108 6 data_in[185]
port 98 nsew signal input
rlabel metal2 s 54574 78308 54630 79108 6 data_in[186]
port 99 nsew signal input
rlabel metal2 s 54850 78308 54906 79108 6 data_in[187]
port 100 nsew signal input
rlabel metal2 s 55126 78308 55182 79108 6 data_in[188]
port 101 nsew signal input
rlabel metal2 s 55402 78308 55458 79108 6 data_in[189]
port 102 nsew signal input
rlabel metal2 s 8206 78308 8262 79108 6 data_in[18]
port 103 nsew signal input
rlabel metal2 s 55678 78308 55734 79108 6 data_in[190]
port 104 nsew signal input
rlabel metal2 s 55954 78308 56010 79108 6 data_in[191]
port 105 nsew signal input
rlabel metal2 s 56230 78308 56286 79108 6 data_in[192]
port 106 nsew signal input
rlabel metal2 s 56506 78308 56562 79108 6 data_in[193]
port 107 nsew signal input
rlabel metal2 s 56782 78308 56838 79108 6 data_in[194]
port 108 nsew signal input
rlabel metal2 s 57058 78308 57114 79108 6 data_in[195]
port 109 nsew signal input
rlabel metal2 s 57334 78308 57390 79108 6 data_in[196]
port 110 nsew signal input
rlabel metal2 s 57610 78308 57666 79108 6 data_in[197]
port 111 nsew signal input
rlabel metal2 s 57886 78308 57942 79108 6 data_in[198]
port 112 nsew signal input
rlabel metal2 s 58162 78308 58218 79108 6 data_in[199]
port 113 nsew signal input
rlabel metal2 s 8482 78308 8538 79108 6 data_in[19]
port 114 nsew signal input
rlabel metal2 s 3514 78308 3570 79108 6 data_in[1]
port 115 nsew signal input
rlabel metal2 s 58438 78308 58494 79108 6 data_in[200]
port 116 nsew signal input
rlabel metal2 s 58714 78308 58770 79108 6 data_in[201]
port 117 nsew signal input
rlabel metal2 s 58990 78308 59046 79108 6 data_in[202]
port 118 nsew signal input
rlabel metal2 s 59266 78308 59322 79108 6 data_in[203]
port 119 nsew signal input
rlabel metal2 s 59542 78308 59598 79108 6 data_in[204]
port 120 nsew signal input
rlabel metal2 s 59818 78308 59874 79108 6 data_in[205]
port 121 nsew signal input
rlabel metal2 s 60094 78308 60150 79108 6 data_in[206]
port 122 nsew signal input
rlabel metal2 s 60370 78308 60426 79108 6 data_in[207]
port 123 nsew signal input
rlabel metal2 s 60646 78308 60702 79108 6 data_in[208]
port 124 nsew signal input
rlabel metal2 s 60922 78308 60978 79108 6 data_in[209]
port 125 nsew signal input
rlabel metal2 s 8758 78308 8814 79108 6 data_in[20]
port 126 nsew signal input
rlabel metal2 s 61198 78308 61254 79108 6 data_in[210]
port 127 nsew signal input
rlabel metal2 s 61474 78308 61530 79108 6 data_in[211]
port 128 nsew signal input
rlabel metal2 s 61750 78308 61806 79108 6 data_in[212]
port 129 nsew signal input
rlabel metal2 s 62026 78308 62082 79108 6 data_in[213]
port 130 nsew signal input
rlabel metal2 s 62302 78308 62358 79108 6 data_in[214]
port 131 nsew signal input
rlabel metal2 s 62578 78308 62634 79108 6 data_in[215]
port 132 nsew signal input
rlabel metal2 s 62854 78308 62910 79108 6 data_in[216]
port 133 nsew signal input
rlabel metal2 s 63130 78308 63186 79108 6 data_in[217]
port 134 nsew signal input
rlabel metal2 s 63406 78308 63462 79108 6 data_in[218]
port 135 nsew signal input
rlabel metal2 s 63682 78308 63738 79108 6 data_in[219]
port 136 nsew signal input
rlabel metal2 s 9034 78308 9090 79108 6 data_in[21]
port 137 nsew signal input
rlabel metal2 s 63958 78308 64014 79108 6 data_in[220]
port 138 nsew signal input
rlabel metal2 s 64234 78308 64290 79108 6 data_in[221]
port 139 nsew signal input
rlabel metal2 s 64510 78308 64566 79108 6 data_in[222]
port 140 nsew signal input
rlabel metal2 s 64786 78308 64842 79108 6 data_in[223]
port 141 nsew signal input
rlabel metal2 s 65062 78308 65118 79108 6 data_in[224]
port 142 nsew signal input
rlabel metal2 s 65338 78308 65394 79108 6 data_in[225]
port 143 nsew signal input
rlabel metal2 s 65614 78308 65670 79108 6 data_in[226]
port 144 nsew signal input
rlabel metal2 s 65890 78308 65946 79108 6 data_in[227]
port 145 nsew signal input
rlabel metal2 s 66166 78308 66222 79108 6 data_in[228]
port 146 nsew signal input
rlabel metal2 s 66442 78308 66498 79108 6 data_in[229]
port 147 nsew signal input
rlabel metal2 s 9310 78308 9366 79108 6 data_in[22]
port 148 nsew signal input
rlabel metal2 s 66718 78308 66774 79108 6 data_in[230]
port 149 nsew signal input
rlabel metal2 s 66994 78308 67050 79108 6 data_in[231]
port 150 nsew signal input
rlabel metal2 s 67270 78308 67326 79108 6 data_in[232]
port 151 nsew signal input
rlabel metal2 s 67546 78308 67602 79108 6 data_in[233]
port 152 nsew signal input
rlabel metal2 s 67822 78308 67878 79108 6 data_in[234]
port 153 nsew signal input
rlabel metal2 s 68098 78308 68154 79108 6 data_in[235]
port 154 nsew signal input
rlabel metal2 s 68374 78308 68430 79108 6 data_in[236]
port 155 nsew signal input
rlabel metal2 s 68650 78308 68706 79108 6 data_in[237]
port 156 nsew signal input
rlabel metal2 s 68926 78308 68982 79108 6 data_in[238]
port 157 nsew signal input
rlabel metal2 s 69202 78308 69258 79108 6 data_in[239]
port 158 nsew signal input
rlabel metal2 s 9586 78308 9642 79108 6 data_in[23]
port 159 nsew signal input
rlabel metal2 s 69478 78308 69534 79108 6 data_in[240]
port 160 nsew signal input
rlabel metal2 s 69754 78308 69810 79108 6 data_in[241]
port 161 nsew signal input
rlabel metal2 s 70030 78308 70086 79108 6 data_in[242]
port 162 nsew signal input
rlabel metal2 s 70306 78308 70362 79108 6 data_in[243]
port 163 nsew signal input
rlabel metal2 s 70582 78308 70638 79108 6 data_in[244]
port 164 nsew signal input
rlabel metal2 s 70858 78308 70914 79108 6 data_in[245]
port 165 nsew signal input
rlabel metal2 s 71134 78308 71190 79108 6 data_in[246]
port 166 nsew signal input
rlabel metal2 s 71410 78308 71466 79108 6 data_in[247]
port 167 nsew signal input
rlabel metal2 s 71686 78308 71742 79108 6 data_in[248]
port 168 nsew signal input
rlabel metal2 s 71962 78308 72018 79108 6 data_in[249]
port 169 nsew signal input
rlabel metal2 s 9862 78308 9918 79108 6 data_in[24]
port 170 nsew signal input
rlabel metal2 s 72238 78308 72294 79108 6 data_in[250]
port 171 nsew signal input
rlabel metal2 s 72514 78308 72570 79108 6 data_in[251]
port 172 nsew signal input
rlabel metal2 s 72790 78308 72846 79108 6 data_in[252]
port 173 nsew signal input
rlabel metal2 s 73066 78308 73122 79108 6 data_in[253]
port 174 nsew signal input
rlabel metal2 s 73342 78308 73398 79108 6 data_in[254]
port 175 nsew signal input
rlabel metal2 s 73618 78308 73674 79108 6 data_in[255]
port 176 nsew signal input
rlabel metal2 s 10138 78308 10194 79108 6 data_in[25]
port 177 nsew signal input
rlabel metal2 s 10414 78308 10470 79108 6 data_in[26]
port 178 nsew signal input
rlabel metal2 s 10690 78308 10746 79108 6 data_in[27]
port 179 nsew signal input
rlabel metal2 s 10966 78308 11022 79108 6 data_in[28]
port 180 nsew signal input
rlabel metal2 s 11242 78308 11298 79108 6 data_in[29]
port 181 nsew signal input
rlabel metal2 s 3790 78308 3846 79108 6 data_in[2]
port 182 nsew signal input
rlabel metal2 s 11518 78308 11574 79108 6 data_in[30]
port 183 nsew signal input
rlabel metal2 s 11794 78308 11850 79108 6 data_in[31]
port 184 nsew signal input
rlabel metal2 s 12070 78308 12126 79108 6 data_in[32]
port 185 nsew signal input
rlabel metal2 s 12346 78308 12402 79108 6 data_in[33]
port 186 nsew signal input
rlabel metal2 s 12622 78308 12678 79108 6 data_in[34]
port 187 nsew signal input
rlabel metal2 s 12898 78308 12954 79108 6 data_in[35]
port 188 nsew signal input
rlabel metal2 s 13174 78308 13230 79108 6 data_in[36]
port 189 nsew signal input
rlabel metal2 s 13450 78308 13506 79108 6 data_in[37]
port 190 nsew signal input
rlabel metal2 s 13726 78308 13782 79108 6 data_in[38]
port 191 nsew signal input
rlabel metal2 s 14002 78308 14058 79108 6 data_in[39]
port 192 nsew signal input
rlabel metal2 s 4066 78308 4122 79108 6 data_in[3]
port 193 nsew signal input
rlabel metal2 s 14278 78308 14334 79108 6 data_in[40]
port 194 nsew signal input
rlabel metal2 s 14554 78308 14610 79108 6 data_in[41]
port 195 nsew signal input
rlabel metal2 s 14830 78308 14886 79108 6 data_in[42]
port 196 nsew signal input
rlabel metal2 s 15106 78308 15162 79108 6 data_in[43]
port 197 nsew signal input
rlabel metal2 s 15382 78308 15438 79108 6 data_in[44]
port 198 nsew signal input
rlabel metal2 s 15658 78308 15714 79108 6 data_in[45]
port 199 nsew signal input
rlabel metal2 s 15934 78308 15990 79108 6 data_in[46]
port 200 nsew signal input
rlabel metal2 s 16210 78308 16266 79108 6 data_in[47]
port 201 nsew signal input
rlabel metal2 s 16486 78308 16542 79108 6 data_in[48]
port 202 nsew signal input
rlabel metal2 s 16762 78308 16818 79108 6 data_in[49]
port 203 nsew signal input
rlabel metal2 s 4342 78308 4398 79108 6 data_in[4]
port 204 nsew signal input
rlabel metal2 s 17038 78308 17094 79108 6 data_in[50]
port 205 nsew signal input
rlabel metal2 s 17314 78308 17370 79108 6 data_in[51]
port 206 nsew signal input
rlabel metal2 s 17590 78308 17646 79108 6 data_in[52]
port 207 nsew signal input
rlabel metal2 s 17866 78308 17922 79108 6 data_in[53]
port 208 nsew signal input
rlabel metal2 s 18142 78308 18198 79108 6 data_in[54]
port 209 nsew signal input
rlabel metal2 s 18418 78308 18474 79108 6 data_in[55]
port 210 nsew signal input
rlabel metal2 s 18694 78308 18750 79108 6 data_in[56]
port 211 nsew signal input
rlabel metal2 s 18970 78308 19026 79108 6 data_in[57]
port 212 nsew signal input
rlabel metal2 s 19246 78308 19302 79108 6 data_in[58]
port 213 nsew signal input
rlabel metal2 s 19522 78308 19578 79108 6 data_in[59]
port 214 nsew signal input
rlabel metal2 s 4618 78308 4674 79108 6 data_in[5]
port 215 nsew signal input
rlabel metal2 s 19798 78308 19854 79108 6 data_in[60]
port 216 nsew signal input
rlabel metal2 s 20074 78308 20130 79108 6 data_in[61]
port 217 nsew signal input
rlabel metal2 s 20350 78308 20406 79108 6 data_in[62]
port 218 nsew signal input
rlabel metal2 s 20626 78308 20682 79108 6 data_in[63]
port 219 nsew signal input
rlabel metal2 s 20902 78308 20958 79108 6 data_in[64]
port 220 nsew signal input
rlabel metal2 s 21178 78308 21234 79108 6 data_in[65]
port 221 nsew signal input
rlabel metal2 s 21454 78308 21510 79108 6 data_in[66]
port 222 nsew signal input
rlabel metal2 s 21730 78308 21786 79108 6 data_in[67]
port 223 nsew signal input
rlabel metal2 s 22006 78308 22062 79108 6 data_in[68]
port 224 nsew signal input
rlabel metal2 s 22282 78308 22338 79108 6 data_in[69]
port 225 nsew signal input
rlabel metal2 s 4894 78308 4950 79108 6 data_in[6]
port 226 nsew signal input
rlabel metal2 s 22558 78308 22614 79108 6 data_in[70]
port 227 nsew signal input
rlabel metal2 s 22834 78308 22890 79108 6 data_in[71]
port 228 nsew signal input
rlabel metal2 s 23110 78308 23166 79108 6 data_in[72]
port 229 nsew signal input
rlabel metal2 s 23386 78308 23442 79108 6 data_in[73]
port 230 nsew signal input
rlabel metal2 s 23662 78308 23718 79108 6 data_in[74]
port 231 nsew signal input
rlabel metal2 s 23938 78308 23994 79108 6 data_in[75]
port 232 nsew signal input
rlabel metal2 s 24214 78308 24270 79108 6 data_in[76]
port 233 nsew signal input
rlabel metal2 s 24490 78308 24546 79108 6 data_in[77]
port 234 nsew signal input
rlabel metal2 s 24766 78308 24822 79108 6 data_in[78]
port 235 nsew signal input
rlabel metal2 s 25042 78308 25098 79108 6 data_in[79]
port 236 nsew signal input
rlabel metal2 s 5170 78308 5226 79108 6 data_in[7]
port 237 nsew signal input
rlabel metal2 s 25318 78308 25374 79108 6 data_in[80]
port 238 nsew signal input
rlabel metal2 s 25594 78308 25650 79108 6 data_in[81]
port 239 nsew signal input
rlabel metal2 s 25870 78308 25926 79108 6 data_in[82]
port 240 nsew signal input
rlabel metal2 s 26146 78308 26202 79108 6 data_in[83]
port 241 nsew signal input
rlabel metal2 s 26422 78308 26478 79108 6 data_in[84]
port 242 nsew signal input
rlabel metal2 s 26698 78308 26754 79108 6 data_in[85]
port 243 nsew signal input
rlabel metal2 s 26974 78308 27030 79108 6 data_in[86]
port 244 nsew signal input
rlabel metal2 s 27250 78308 27306 79108 6 data_in[87]
port 245 nsew signal input
rlabel metal2 s 27526 78308 27582 79108 6 data_in[88]
port 246 nsew signal input
rlabel metal2 s 27802 78308 27858 79108 6 data_in[89]
port 247 nsew signal input
rlabel metal2 s 5446 78308 5502 79108 6 data_in[8]
port 248 nsew signal input
rlabel metal2 s 28078 78308 28134 79108 6 data_in[90]
port 249 nsew signal input
rlabel metal2 s 28354 78308 28410 79108 6 data_in[91]
port 250 nsew signal input
rlabel metal2 s 28630 78308 28686 79108 6 data_in[92]
port 251 nsew signal input
rlabel metal2 s 28906 78308 28962 79108 6 data_in[93]
port 252 nsew signal input
rlabel metal2 s 29182 78308 29238 79108 6 data_in[94]
port 253 nsew signal input
rlabel metal2 s 29458 78308 29514 79108 6 data_in[95]
port 254 nsew signal input
rlabel metal2 s 29734 78308 29790 79108 6 data_in[96]
port 255 nsew signal input
rlabel metal2 s 30010 78308 30066 79108 6 data_in[97]
port 256 nsew signal input
rlabel metal2 s 30286 78308 30342 79108 6 data_in[98]
port 257 nsew signal input
rlabel metal2 s 30562 78308 30618 79108 6 data_in[99]
port 258 nsew signal input
rlabel metal2 s 5722 78308 5778 79108 6 data_in[9]
port 259 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 data_out[0]
port 260 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 data_out[10]
port 261 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 data_out[11]
port 262 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 data_out[12]
port 263 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 data_out[13]
port 264 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 data_out[14]
port 265 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 data_out[15]
port 266 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 data_out[16]
port 267 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 data_out[17]
port 268 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 data_out[18]
port 269 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 data_out[19]
port 270 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 data_out[1]
port 271 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 data_out[20]
port 272 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 data_out[21]
port 273 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 data_out[22]
port 274 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 data_out[23]
port 275 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 data_out[24]
port 276 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 data_out[25]
port 277 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 data_out[26]
port 278 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 data_out[27]
port 279 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 data_out[2]
port 280 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 data_out[3]
port 281 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 data_out[4]
port 282 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 data_out[5]
port 283 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 data_out[6]
port 284 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 data_out[7]
port 285 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 data_out[8]
port 286 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 data_out[9]
port 287 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 reset
port 288 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 76964 79108
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17635744
string GDS_FILE /home/ucass/Work/DNN_ACC_IITGN/openlane/mac/runs/23_09_22_02_42/results/signoff/mac.magic.gds
string GDS_START 1055784
<< end >>

