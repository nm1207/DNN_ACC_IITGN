magic
tech sky130A
magscale 1 2
timestamp 1695414633
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 212 558978 349840
<< metal2 >>
rect 7838 0 7894 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17774 0 17830 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28814 0 28870 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32126 0 32182 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47582 0 47638 800
rect 48686 0 48742 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56414 0 56470 800
rect 57518 0 57574 800
rect 58622 0 58678 800
rect 59726 0 59782 800
rect 60830 0 60886 800
rect 61934 0 61990 800
rect 63038 0 63094 800
rect 64142 0 64198 800
rect 65246 0 65302 800
rect 66350 0 66406 800
rect 67454 0 67510 800
rect 68558 0 68614 800
rect 69662 0 69718 800
rect 70766 0 70822 800
rect 71870 0 71926 800
rect 72974 0 73030 800
rect 74078 0 74134 800
rect 75182 0 75238 800
rect 76286 0 76342 800
rect 77390 0 77446 800
rect 78494 0 78550 800
rect 79598 0 79654 800
rect 80702 0 80758 800
rect 81806 0 81862 800
rect 82910 0 82966 800
rect 84014 0 84070 800
rect 85118 0 85174 800
rect 86222 0 86278 800
rect 87326 0 87382 800
rect 88430 0 88486 800
rect 89534 0 89590 800
rect 90638 0 90694 800
rect 91742 0 91798 800
rect 92846 0 92902 800
rect 93950 0 94006 800
rect 95054 0 95110 800
rect 96158 0 96214 800
rect 97262 0 97318 800
rect 98366 0 98422 800
rect 99470 0 99526 800
rect 100574 0 100630 800
rect 101678 0 101734 800
rect 102782 0 102838 800
rect 103886 0 103942 800
rect 104990 0 105046 800
rect 106094 0 106150 800
rect 107198 0 107254 800
rect 108302 0 108358 800
rect 109406 0 109462 800
rect 110510 0 110566 800
rect 111614 0 111670 800
rect 112718 0 112774 800
rect 113822 0 113878 800
rect 114926 0 114982 800
rect 116030 0 116086 800
rect 117134 0 117190 800
rect 118238 0 118294 800
rect 119342 0 119398 800
rect 120446 0 120502 800
rect 121550 0 121606 800
rect 122654 0 122710 800
rect 123758 0 123814 800
rect 124862 0 124918 800
rect 125966 0 126022 800
rect 127070 0 127126 800
rect 128174 0 128230 800
rect 129278 0 129334 800
rect 130382 0 130438 800
rect 131486 0 131542 800
rect 132590 0 132646 800
rect 133694 0 133750 800
rect 134798 0 134854 800
rect 135902 0 135958 800
rect 137006 0 137062 800
rect 138110 0 138166 800
rect 139214 0 139270 800
rect 140318 0 140374 800
rect 141422 0 141478 800
rect 142526 0 142582 800
rect 143630 0 143686 800
rect 144734 0 144790 800
rect 145838 0 145894 800
rect 146942 0 146998 800
rect 148046 0 148102 800
rect 149150 0 149206 800
rect 150254 0 150310 800
rect 151358 0 151414 800
rect 152462 0 152518 800
rect 153566 0 153622 800
rect 154670 0 154726 800
rect 155774 0 155830 800
rect 156878 0 156934 800
rect 157982 0 158038 800
rect 159086 0 159142 800
rect 160190 0 160246 800
rect 161294 0 161350 800
rect 162398 0 162454 800
rect 163502 0 163558 800
rect 164606 0 164662 800
rect 165710 0 165766 800
rect 166814 0 166870 800
rect 167918 0 167974 800
rect 169022 0 169078 800
rect 170126 0 170182 800
rect 171230 0 171286 800
rect 172334 0 172390 800
rect 173438 0 173494 800
rect 174542 0 174598 800
rect 175646 0 175702 800
rect 176750 0 176806 800
rect 177854 0 177910 800
rect 178958 0 179014 800
rect 180062 0 180118 800
rect 181166 0 181222 800
rect 182270 0 182326 800
rect 183374 0 183430 800
rect 184478 0 184534 800
rect 185582 0 185638 800
rect 186686 0 186742 800
rect 187790 0 187846 800
rect 188894 0 188950 800
rect 189998 0 190054 800
rect 191102 0 191158 800
rect 192206 0 192262 800
rect 193310 0 193366 800
rect 194414 0 194470 800
rect 195518 0 195574 800
rect 196622 0 196678 800
rect 197726 0 197782 800
rect 198830 0 198886 800
rect 199934 0 199990 800
rect 201038 0 201094 800
rect 202142 0 202198 800
rect 203246 0 203302 800
rect 204350 0 204406 800
rect 205454 0 205510 800
rect 206558 0 206614 800
rect 207662 0 207718 800
rect 208766 0 208822 800
rect 209870 0 209926 800
rect 210974 0 211030 800
rect 212078 0 212134 800
rect 213182 0 213238 800
rect 214286 0 214342 800
rect 215390 0 215446 800
rect 216494 0 216550 800
rect 217598 0 217654 800
rect 218702 0 218758 800
rect 219806 0 219862 800
rect 220910 0 220966 800
rect 222014 0 222070 800
rect 223118 0 223174 800
rect 224222 0 224278 800
rect 225326 0 225382 800
rect 226430 0 226486 800
rect 227534 0 227590 800
rect 228638 0 228694 800
rect 229742 0 229798 800
rect 230846 0 230902 800
rect 231950 0 232006 800
rect 233054 0 233110 800
rect 234158 0 234214 800
rect 235262 0 235318 800
rect 236366 0 236422 800
rect 237470 0 237526 800
rect 238574 0 238630 800
rect 239678 0 239734 800
rect 240782 0 240838 800
rect 241886 0 241942 800
rect 242990 0 243046 800
rect 244094 0 244150 800
rect 245198 0 245254 800
rect 246302 0 246358 800
rect 247406 0 247462 800
rect 248510 0 248566 800
rect 249614 0 249670 800
rect 250718 0 250774 800
rect 251822 0 251878 800
rect 252926 0 252982 800
rect 254030 0 254086 800
rect 255134 0 255190 800
rect 256238 0 256294 800
rect 257342 0 257398 800
rect 258446 0 258502 800
rect 259550 0 259606 800
rect 260654 0 260710 800
rect 261758 0 261814 800
rect 262862 0 262918 800
rect 263966 0 264022 800
rect 265070 0 265126 800
rect 266174 0 266230 800
rect 267278 0 267334 800
rect 268382 0 268438 800
rect 269486 0 269542 800
rect 270590 0 270646 800
rect 271694 0 271750 800
rect 272798 0 272854 800
rect 273902 0 273958 800
rect 275006 0 275062 800
rect 276110 0 276166 800
rect 277214 0 277270 800
rect 278318 0 278374 800
rect 279422 0 279478 800
rect 280526 0 280582 800
rect 281630 0 281686 800
rect 282734 0 282790 800
rect 283838 0 283894 800
rect 284942 0 284998 800
rect 286046 0 286102 800
rect 287150 0 287206 800
rect 288254 0 288310 800
rect 289358 0 289414 800
rect 290462 0 290518 800
rect 291566 0 291622 800
rect 292670 0 292726 800
rect 293774 0 293830 800
rect 294878 0 294934 800
rect 295982 0 296038 800
rect 297086 0 297142 800
rect 298190 0 298246 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301502 0 301558 800
rect 302606 0 302662 800
rect 303710 0 303766 800
rect 304814 0 304870 800
rect 305918 0 305974 800
rect 307022 0 307078 800
rect 308126 0 308182 800
rect 309230 0 309286 800
rect 310334 0 310390 800
rect 311438 0 311494 800
rect 312542 0 312598 800
rect 313646 0 313702 800
rect 314750 0 314806 800
rect 315854 0 315910 800
rect 316958 0 317014 800
rect 318062 0 318118 800
rect 319166 0 319222 800
rect 320270 0 320326 800
rect 321374 0 321430 800
rect 322478 0 322534 800
rect 323582 0 323638 800
rect 324686 0 324742 800
rect 325790 0 325846 800
rect 326894 0 326950 800
rect 327998 0 328054 800
rect 329102 0 329158 800
rect 330206 0 330262 800
rect 331310 0 331366 800
rect 332414 0 332470 800
rect 333518 0 333574 800
rect 334622 0 334678 800
rect 335726 0 335782 800
rect 336830 0 336886 800
rect 337934 0 337990 800
rect 339038 0 339094 800
rect 340142 0 340198 800
rect 341246 0 341302 800
rect 342350 0 342406 800
rect 343454 0 343510 800
rect 344558 0 344614 800
rect 345662 0 345718 800
rect 346766 0 346822 800
rect 347870 0 347926 800
rect 348974 0 349030 800
rect 350078 0 350134 800
rect 351182 0 351238 800
rect 352286 0 352342 800
rect 353390 0 353446 800
rect 354494 0 354550 800
rect 355598 0 355654 800
rect 356702 0 356758 800
rect 357806 0 357862 800
rect 358910 0 358966 800
rect 360014 0 360070 800
rect 361118 0 361174 800
rect 362222 0 362278 800
rect 363326 0 363382 800
rect 364430 0 364486 800
rect 365534 0 365590 800
rect 366638 0 366694 800
rect 367742 0 367798 800
rect 368846 0 368902 800
rect 369950 0 370006 800
rect 371054 0 371110 800
rect 372158 0 372214 800
rect 373262 0 373318 800
rect 374366 0 374422 800
rect 375470 0 375526 800
rect 376574 0 376630 800
rect 377678 0 377734 800
rect 378782 0 378838 800
rect 379886 0 379942 800
rect 380990 0 381046 800
rect 382094 0 382150 800
rect 383198 0 383254 800
rect 384302 0 384358 800
rect 385406 0 385462 800
rect 386510 0 386566 800
rect 387614 0 387670 800
rect 388718 0 388774 800
rect 389822 0 389878 800
rect 390926 0 390982 800
rect 392030 0 392086 800
rect 393134 0 393190 800
rect 394238 0 394294 800
rect 395342 0 395398 800
rect 396446 0 396502 800
rect 397550 0 397606 800
rect 398654 0 398710 800
rect 399758 0 399814 800
rect 400862 0 400918 800
rect 401966 0 402022 800
rect 403070 0 403126 800
rect 404174 0 404230 800
rect 405278 0 405334 800
rect 406382 0 406438 800
rect 407486 0 407542 800
rect 408590 0 408646 800
rect 409694 0 409750 800
rect 410798 0 410854 800
rect 411902 0 411958 800
rect 413006 0 413062 800
rect 414110 0 414166 800
rect 415214 0 415270 800
rect 416318 0 416374 800
rect 417422 0 417478 800
rect 418526 0 418582 800
rect 419630 0 419686 800
rect 420734 0 420790 800
rect 421838 0 421894 800
rect 422942 0 422998 800
rect 424046 0 424102 800
rect 425150 0 425206 800
rect 426254 0 426310 800
rect 427358 0 427414 800
rect 428462 0 428518 800
rect 429566 0 429622 800
rect 430670 0 430726 800
rect 431774 0 431830 800
rect 432878 0 432934 800
rect 433982 0 434038 800
rect 435086 0 435142 800
rect 436190 0 436246 800
rect 437294 0 437350 800
rect 438398 0 438454 800
rect 439502 0 439558 800
rect 440606 0 440662 800
rect 441710 0 441766 800
rect 442814 0 442870 800
rect 443918 0 443974 800
rect 445022 0 445078 800
rect 446126 0 446182 800
rect 447230 0 447286 800
rect 448334 0 448390 800
rect 449438 0 449494 800
rect 450542 0 450598 800
rect 451646 0 451702 800
rect 452750 0 452806 800
rect 453854 0 453910 800
rect 454958 0 455014 800
rect 456062 0 456118 800
rect 457166 0 457222 800
rect 458270 0 458326 800
rect 459374 0 459430 800
rect 460478 0 460534 800
rect 461582 0 461638 800
rect 462686 0 462742 800
rect 463790 0 463846 800
rect 464894 0 464950 800
rect 465998 0 466054 800
rect 467102 0 467158 800
rect 468206 0 468262 800
rect 469310 0 469366 800
rect 470414 0 470470 800
rect 471518 0 471574 800
rect 472622 0 472678 800
rect 473726 0 473782 800
rect 474830 0 474886 800
rect 475934 0 475990 800
rect 477038 0 477094 800
rect 478142 0 478198 800
rect 479246 0 479302 800
rect 480350 0 480406 800
rect 481454 0 481510 800
rect 482558 0 482614 800
rect 483662 0 483718 800
rect 484766 0 484822 800
rect 485870 0 485926 800
rect 486974 0 487030 800
rect 488078 0 488134 800
rect 489182 0 489238 800
rect 490286 0 490342 800
rect 491390 0 491446 800
rect 492494 0 492550 800
rect 493598 0 493654 800
rect 494702 0 494758 800
rect 495806 0 495862 800
rect 496910 0 496966 800
rect 498014 0 498070 800
rect 499118 0 499174 800
rect 500222 0 500278 800
rect 501326 0 501382 800
rect 502430 0 502486 800
rect 503534 0 503590 800
rect 504638 0 504694 800
rect 505742 0 505798 800
rect 506846 0 506902 800
rect 507950 0 508006 800
rect 509054 0 509110 800
rect 510158 0 510214 800
rect 511262 0 511318 800
rect 512366 0 512422 800
rect 513470 0 513526 800
rect 514574 0 514630 800
rect 515678 0 515734 800
rect 516782 0 516838 800
rect 517886 0 517942 800
rect 518990 0 519046 800
rect 520094 0 520150 800
rect 521198 0 521254 800
rect 522302 0 522358 800
rect 523406 0 523462 800
rect 524510 0 524566 800
rect 525614 0 525670 800
rect 526718 0 526774 800
rect 527822 0 527878 800
rect 528926 0 528982 800
rect 530030 0 530086 800
rect 531134 0 531190 800
rect 532238 0 532294 800
rect 533342 0 533398 800
rect 534446 0 534502 800
rect 535550 0 535606 800
rect 536654 0 536710 800
rect 537758 0 537814 800
rect 538862 0 538918 800
rect 539966 0 540022 800
rect 541070 0 541126 800
rect 542174 0 542230 800
rect 543278 0 543334 800
rect 544382 0 544438 800
rect 545486 0 545542 800
rect 546590 0 546646 800
rect 547694 0 547750 800
rect 548798 0 548854 800
rect 549902 0 549958 800
rect 551006 0 551062 800
rect 552110 0 552166 800
<< obsm2 >>
rect 938 856 558974 349829
rect 938 167 7782 856
rect 7950 167 8886 856
rect 9054 167 9990 856
rect 10158 167 11094 856
rect 11262 167 12198 856
rect 12366 167 13302 856
rect 13470 167 14406 856
rect 14574 167 15510 856
rect 15678 167 16614 856
rect 16782 167 17718 856
rect 17886 167 18822 856
rect 18990 167 19926 856
rect 20094 167 21030 856
rect 21198 167 22134 856
rect 22302 167 23238 856
rect 23406 167 24342 856
rect 24510 167 25446 856
rect 25614 167 26550 856
rect 26718 167 27654 856
rect 27822 167 28758 856
rect 28926 167 29862 856
rect 30030 167 30966 856
rect 31134 167 32070 856
rect 32238 167 33174 856
rect 33342 167 34278 856
rect 34446 167 35382 856
rect 35550 167 36486 856
rect 36654 167 37590 856
rect 37758 167 38694 856
rect 38862 167 39798 856
rect 39966 167 40902 856
rect 41070 167 42006 856
rect 42174 167 43110 856
rect 43278 167 44214 856
rect 44382 167 45318 856
rect 45486 167 46422 856
rect 46590 167 47526 856
rect 47694 167 48630 856
rect 48798 167 49734 856
rect 49902 167 50838 856
rect 51006 167 51942 856
rect 52110 167 53046 856
rect 53214 167 54150 856
rect 54318 167 55254 856
rect 55422 167 56358 856
rect 56526 167 57462 856
rect 57630 167 58566 856
rect 58734 167 59670 856
rect 59838 167 60774 856
rect 60942 167 61878 856
rect 62046 167 62982 856
rect 63150 167 64086 856
rect 64254 167 65190 856
rect 65358 167 66294 856
rect 66462 167 67398 856
rect 67566 167 68502 856
rect 68670 167 69606 856
rect 69774 167 70710 856
rect 70878 167 71814 856
rect 71982 167 72918 856
rect 73086 167 74022 856
rect 74190 167 75126 856
rect 75294 167 76230 856
rect 76398 167 77334 856
rect 77502 167 78438 856
rect 78606 167 79542 856
rect 79710 167 80646 856
rect 80814 167 81750 856
rect 81918 167 82854 856
rect 83022 167 83958 856
rect 84126 167 85062 856
rect 85230 167 86166 856
rect 86334 167 87270 856
rect 87438 167 88374 856
rect 88542 167 89478 856
rect 89646 167 90582 856
rect 90750 167 91686 856
rect 91854 167 92790 856
rect 92958 167 93894 856
rect 94062 167 94998 856
rect 95166 167 96102 856
rect 96270 167 97206 856
rect 97374 167 98310 856
rect 98478 167 99414 856
rect 99582 167 100518 856
rect 100686 167 101622 856
rect 101790 167 102726 856
rect 102894 167 103830 856
rect 103998 167 104934 856
rect 105102 167 106038 856
rect 106206 167 107142 856
rect 107310 167 108246 856
rect 108414 167 109350 856
rect 109518 167 110454 856
rect 110622 167 111558 856
rect 111726 167 112662 856
rect 112830 167 113766 856
rect 113934 167 114870 856
rect 115038 167 115974 856
rect 116142 167 117078 856
rect 117246 167 118182 856
rect 118350 167 119286 856
rect 119454 167 120390 856
rect 120558 167 121494 856
rect 121662 167 122598 856
rect 122766 167 123702 856
rect 123870 167 124806 856
rect 124974 167 125910 856
rect 126078 167 127014 856
rect 127182 167 128118 856
rect 128286 167 129222 856
rect 129390 167 130326 856
rect 130494 167 131430 856
rect 131598 167 132534 856
rect 132702 167 133638 856
rect 133806 167 134742 856
rect 134910 167 135846 856
rect 136014 167 136950 856
rect 137118 167 138054 856
rect 138222 167 139158 856
rect 139326 167 140262 856
rect 140430 167 141366 856
rect 141534 167 142470 856
rect 142638 167 143574 856
rect 143742 167 144678 856
rect 144846 167 145782 856
rect 145950 167 146886 856
rect 147054 167 147990 856
rect 148158 167 149094 856
rect 149262 167 150198 856
rect 150366 167 151302 856
rect 151470 167 152406 856
rect 152574 167 153510 856
rect 153678 167 154614 856
rect 154782 167 155718 856
rect 155886 167 156822 856
rect 156990 167 157926 856
rect 158094 167 159030 856
rect 159198 167 160134 856
rect 160302 167 161238 856
rect 161406 167 162342 856
rect 162510 167 163446 856
rect 163614 167 164550 856
rect 164718 167 165654 856
rect 165822 167 166758 856
rect 166926 167 167862 856
rect 168030 167 168966 856
rect 169134 167 170070 856
rect 170238 167 171174 856
rect 171342 167 172278 856
rect 172446 167 173382 856
rect 173550 167 174486 856
rect 174654 167 175590 856
rect 175758 167 176694 856
rect 176862 167 177798 856
rect 177966 167 178902 856
rect 179070 167 180006 856
rect 180174 167 181110 856
rect 181278 167 182214 856
rect 182382 167 183318 856
rect 183486 167 184422 856
rect 184590 167 185526 856
rect 185694 167 186630 856
rect 186798 167 187734 856
rect 187902 167 188838 856
rect 189006 167 189942 856
rect 190110 167 191046 856
rect 191214 167 192150 856
rect 192318 167 193254 856
rect 193422 167 194358 856
rect 194526 167 195462 856
rect 195630 167 196566 856
rect 196734 167 197670 856
rect 197838 167 198774 856
rect 198942 167 199878 856
rect 200046 167 200982 856
rect 201150 167 202086 856
rect 202254 167 203190 856
rect 203358 167 204294 856
rect 204462 167 205398 856
rect 205566 167 206502 856
rect 206670 167 207606 856
rect 207774 167 208710 856
rect 208878 167 209814 856
rect 209982 167 210918 856
rect 211086 167 212022 856
rect 212190 167 213126 856
rect 213294 167 214230 856
rect 214398 167 215334 856
rect 215502 167 216438 856
rect 216606 167 217542 856
rect 217710 167 218646 856
rect 218814 167 219750 856
rect 219918 167 220854 856
rect 221022 167 221958 856
rect 222126 167 223062 856
rect 223230 167 224166 856
rect 224334 167 225270 856
rect 225438 167 226374 856
rect 226542 167 227478 856
rect 227646 167 228582 856
rect 228750 167 229686 856
rect 229854 167 230790 856
rect 230958 167 231894 856
rect 232062 167 232998 856
rect 233166 167 234102 856
rect 234270 167 235206 856
rect 235374 167 236310 856
rect 236478 167 237414 856
rect 237582 167 238518 856
rect 238686 167 239622 856
rect 239790 167 240726 856
rect 240894 167 241830 856
rect 241998 167 242934 856
rect 243102 167 244038 856
rect 244206 167 245142 856
rect 245310 167 246246 856
rect 246414 167 247350 856
rect 247518 167 248454 856
rect 248622 167 249558 856
rect 249726 167 250662 856
rect 250830 167 251766 856
rect 251934 167 252870 856
rect 253038 167 253974 856
rect 254142 167 255078 856
rect 255246 167 256182 856
rect 256350 167 257286 856
rect 257454 167 258390 856
rect 258558 167 259494 856
rect 259662 167 260598 856
rect 260766 167 261702 856
rect 261870 167 262806 856
rect 262974 167 263910 856
rect 264078 167 265014 856
rect 265182 167 266118 856
rect 266286 167 267222 856
rect 267390 167 268326 856
rect 268494 167 269430 856
rect 269598 167 270534 856
rect 270702 167 271638 856
rect 271806 167 272742 856
rect 272910 167 273846 856
rect 274014 167 274950 856
rect 275118 167 276054 856
rect 276222 167 277158 856
rect 277326 167 278262 856
rect 278430 167 279366 856
rect 279534 167 280470 856
rect 280638 167 281574 856
rect 281742 167 282678 856
rect 282846 167 283782 856
rect 283950 167 284886 856
rect 285054 167 285990 856
rect 286158 167 287094 856
rect 287262 167 288198 856
rect 288366 167 289302 856
rect 289470 167 290406 856
rect 290574 167 291510 856
rect 291678 167 292614 856
rect 292782 167 293718 856
rect 293886 167 294822 856
rect 294990 167 295926 856
rect 296094 167 297030 856
rect 297198 167 298134 856
rect 298302 167 299238 856
rect 299406 167 300342 856
rect 300510 167 301446 856
rect 301614 167 302550 856
rect 302718 167 303654 856
rect 303822 167 304758 856
rect 304926 167 305862 856
rect 306030 167 306966 856
rect 307134 167 308070 856
rect 308238 167 309174 856
rect 309342 167 310278 856
rect 310446 167 311382 856
rect 311550 167 312486 856
rect 312654 167 313590 856
rect 313758 167 314694 856
rect 314862 167 315798 856
rect 315966 167 316902 856
rect 317070 167 318006 856
rect 318174 167 319110 856
rect 319278 167 320214 856
rect 320382 167 321318 856
rect 321486 167 322422 856
rect 322590 167 323526 856
rect 323694 167 324630 856
rect 324798 167 325734 856
rect 325902 167 326838 856
rect 327006 167 327942 856
rect 328110 167 329046 856
rect 329214 167 330150 856
rect 330318 167 331254 856
rect 331422 167 332358 856
rect 332526 167 333462 856
rect 333630 167 334566 856
rect 334734 167 335670 856
rect 335838 167 336774 856
rect 336942 167 337878 856
rect 338046 167 338982 856
rect 339150 167 340086 856
rect 340254 167 341190 856
rect 341358 167 342294 856
rect 342462 167 343398 856
rect 343566 167 344502 856
rect 344670 167 345606 856
rect 345774 167 346710 856
rect 346878 167 347814 856
rect 347982 167 348918 856
rect 349086 167 350022 856
rect 350190 167 351126 856
rect 351294 167 352230 856
rect 352398 167 353334 856
rect 353502 167 354438 856
rect 354606 167 355542 856
rect 355710 167 356646 856
rect 356814 167 357750 856
rect 357918 167 358854 856
rect 359022 167 359958 856
rect 360126 167 361062 856
rect 361230 167 362166 856
rect 362334 167 363270 856
rect 363438 167 364374 856
rect 364542 167 365478 856
rect 365646 167 366582 856
rect 366750 167 367686 856
rect 367854 167 368790 856
rect 368958 167 369894 856
rect 370062 167 370998 856
rect 371166 167 372102 856
rect 372270 167 373206 856
rect 373374 167 374310 856
rect 374478 167 375414 856
rect 375582 167 376518 856
rect 376686 167 377622 856
rect 377790 167 378726 856
rect 378894 167 379830 856
rect 379998 167 380934 856
rect 381102 167 382038 856
rect 382206 167 383142 856
rect 383310 167 384246 856
rect 384414 167 385350 856
rect 385518 167 386454 856
rect 386622 167 387558 856
rect 387726 167 388662 856
rect 388830 167 389766 856
rect 389934 167 390870 856
rect 391038 167 391974 856
rect 392142 167 393078 856
rect 393246 167 394182 856
rect 394350 167 395286 856
rect 395454 167 396390 856
rect 396558 167 397494 856
rect 397662 167 398598 856
rect 398766 167 399702 856
rect 399870 167 400806 856
rect 400974 167 401910 856
rect 402078 167 403014 856
rect 403182 167 404118 856
rect 404286 167 405222 856
rect 405390 167 406326 856
rect 406494 167 407430 856
rect 407598 167 408534 856
rect 408702 167 409638 856
rect 409806 167 410742 856
rect 410910 167 411846 856
rect 412014 167 412950 856
rect 413118 167 414054 856
rect 414222 167 415158 856
rect 415326 167 416262 856
rect 416430 167 417366 856
rect 417534 167 418470 856
rect 418638 167 419574 856
rect 419742 167 420678 856
rect 420846 167 421782 856
rect 421950 167 422886 856
rect 423054 167 423990 856
rect 424158 167 425094 856
rect 425262 167 426198 856
rect 426366 167 427302 856
rect 427470 167 428406 856
rect 428574 167 429510 856
rect 429678 167 430614 856
rect 430782 167 431718 856
rect 431886 167 432822 856
rect 432990 167 433926 856
rect 434094 167 435030 856
rect 435198 167 436134 856
rect 436302 167 437238 856
rect 437406 167 438342 856
rect 438510 167 439446 856
rect 439614 167 440550 856
rect 440718 167 441654 856
rect 441822 167 442758 856
rect 442926 167 443862 856
rect 444030 167 444966 856
rect 445134 167 446070 856
rect 446238 167 447174 856
rect 447342 167 448278 856
rect 448446 167 449382 856
rect 449550 167 450486 856
rect 450654 167 451590 856
rect 451758 167 452694 856
rect 452862 167 453798 856
rect 453966 167 454902 856
rect 455070 167 456006 856
rect 456174 167 457110 856
rect 457278 167 458214 856
rect 458382 167 459318 856
rect 459486 167 460422 856
rect 460590 167 461526 856
rect 461694 167 462630 856
rect 462798 167 463734 856
rect 463902 167 464838 856
rect 465006 167 465942 856
rect 466110 167 467046 856
rect 467214 167 468150 856
rect 468318 167 469254 856
rect 469422 167 470358 856
rect 470526 167 471462 856
rect 471630 167 472566 856
rect 472734 167 473670 856
rect 473838 167 474774 856
rect 474942 167 475878 856
rect 476046 167 476982 856
rect 477150 167 478086 856
rect 478254 167 479190 856
rect 479358 167 480294 856
rect 480462 167 481398 856
rect 481566 167 482502 856
rect 482670 167 483606 856
rect 483774 167 484710 856
rect 484878 167 485814 856
rect 485982 167 486918 856
rect 487086 167 488022 856
rect 488190 167 489126 856
rect 489294 167 490230 856
rect 490398 167 491334 856
rect 491502 167 492438 856
rect 492606 167 493542 856
rect 493710 167 494646 856
rect 494814 167 495750 856
rect 495918 167 496854 856
rect 497022 167 497958 856
rect 498126 167 499062 856
rect 499230 167 500166 856
rect 500334 167 501270 856
rect 501438 167 502374 856
rect 502542 167 503478 856
rect 503646 167 504582 856
rect 504750 167 505686 856
rect 505854 167 506790 856
rect 506958 167 507894 856
rect 508062 167 508998 856
rect 509166 167 510102 856
rect 510270 167 511206 856
rect 511374 167 512310 856
rect 512478 167 513414 856
rect 513582 167 514518 856
rect 514686 167 515622 856
rect 515790 167 516726 856
rect 516894 167 517830 856
rect 517998 167 518934 856
rect 519102 167 520038 856
rect 520206 167 521142 856
rect 521310 167 522246 856
rect 522414 167 523350 856
rect 523518 167 524454 856
rect 524622 167 525558 856
rect 525726 167 526662 856
rect 526830 167 527766 856
rect 527934 167 528870 856
rect 529038 167 529974 856
rect 530142 167 531078 856
rect 531246 167 532182 856
rect 532350 167 533286 856
rect 533454 167 534390 856
rect 534558 167 535494 856
rect 535662 167 536598 856
rect 536766 167 537702 856
rect 537870 167 538806 856
rect 538974 167 539910 856
rect 540078 167 541014 856
rect 541182 167 542118 856
rect 542286 167 543222 856
rect 543390 167 544326 856
rect 544494 167 545430 856
rect 545598 167 546534 856
rect 546702 167 547638 856
rect 547806 167 548742 856
rect 548910 167 549846 856
rect 550014 167 550950 856
rect 551118 167 552054 856
rect 552222 167 558974 856
<< metal3 >>
rect 0 343816 800 343936
rect 559200 341912 560000 342032
rect 0 338648 800 338768
rect 559200 334840 560000 334960
rect 0 333480 800 333600
rect 0 328312 800 328432
rect 559200 327768 560000 327888
rect 0 323144 800 323264
rect 559200 320696 560000 320816
rect 0 317976 800 318096
rect 559200 313624 560000 313744
rect 0 312808 800 312928
rect 0 307640 800 307760
rect 559200 306552 560000 306672
rect 0 302472 800 302592
rect 559200 299480 560000 299600
rect 0 297304 800 297424
rect 559200 292408 560000 292528
rect 0 292136 800 292256
rect 0 286968 800 287088
rect 559200 285336 560000 285456
rect 0 281800 800 281920
rect 559200 278264 560000 278384
rect 0 276632 800 276752
rect 0 271464 800 271584
rect 559200 271192 560000 271312
rect 0 266296 800 266416
rect 559200 264120 560000 264240
rect 0 261128 800 261248
rect 559200 257048 560000 257168
rect 0 255960 800 256080
rect 0 250792 800 250912
rect 559200 249976 560000 250096
rect 0 245624 800 245744
rect 559200 242904 560000 243024
rect 0 240456 800 240576
rect 559200 235832 560000 235952
rect 0 235288 800 235408
rect 0 230120 800 230240
rect 559200 228760 560000 228880
rect 0 224952 800 225072
rect 559200 221688 560000 221808
rect 0 219784 800 219904
rect 0 214616 800 214736
rect 559200 214616 560000 214736
rect 0 209448 800 209568
rect 559200 207544 560000 207664
rect 0 204280 800 204400
rect 559200 200472 560000 200592
rect 0 199112 800 199232
rect 0 193944 800 194064
rect 559200 193400 560000 193520
rect 0 188776 800 188896
rect 559200 186328 560000 186448
rect 0 183608 800 183728
rect 559200 179256 560000 179376
rect 0 178440 800 178560
rect 0 173272 800 173392
rect 559200 172184 560000 172304
rect 0 168104 800 168224
rect 559200 165112 560000 165232
rect 0 162936 800 163056
rect 559200 158040 560000 158160
rect 0 157768 800 157888
rect 0 152600 800 152720
rect 559200 150968 560000 151088
rect 0 147432 800 147552
rect 559200 143896 560000 144016
rect 0 142264 800 142384
rect 0 137096 800 137216
rect 559200 136824 560000 136944
rect 0 131928 800 132048
rect 559200 129752 560000 129872
rect 0 126760 800 126880
rect 559200 122680 560000 122800
rect 0 121592 800 121712
rect 0 116424 800 116544
rect 559200 115608 560000 115728
rect 0 111256 800 111376
rect 559200 108536 560000 108656
rect 0 106088 800 106208
rect 559200 101464 560000 101584
rect 0 100920 800 101040
rect 0 95752 800 95872
rect 559200 94392 560000 94512
rect 0 90584 800 90704
rect 559200 87320 560000 87440
rect 0 85416 800 85536
rect 0 80248 800 80368
rect 559200 80248 560000 80368
rect 0 75080 800 75200
rect 559200 73176 560000 73296
rect 0 69912 800 70032
rect 559200 66104 560000 66224
rect 0 64744 800 64864
rect 0 59576 800 59696
rect 559200 59032 560000 59152
rect 0 54408 800 54528
rect 559200 51960 560000 52080
rect 0 49240 800 49360
rect 559200 44888 560000 45008
rect 0 44072 800 44192
rect 0 38904 800 39024
rect 559200 37816 560000 37936
rect 0 33736 800 33856
rect 559200 30744 560000 30864
rect 0 28568 800 28688
rect 559200 23672 560000 23792
rect 0 23400 800 23520
rect 0 18232 800 18352
rect 559200 16600 560000 16720
rect 0 13064 800 13184
rect 559200 9528 560000 9648
rect 0 7896 800 8016
<< obsm3 >>
rect 798 344016 559200 349825
rect 880 343736 559200 344016
rect 798 342112 559200 343736
rect 798 341832 559120 342112
rect 798 338848 559200 341832
rect 880 338568 559200 338848
rect 798 335040 559200 338568
rect 798 334760 559120 335040
rect 798 333680 559200 334760
rect 880 333400 559200 333680
rect 798 328512 559200 333400
rect 880 328232 559200 328512
rect 798 327968 559200 328232
rect 798 327688 559120 327968
rect 798 323344 559200 327688
rect 880 323064 559200 323344
rect 798 320896 559200 323064
rect 798 320616 559120 320896
rect 798 318176 559200 320616
rect 880 317896 559200 318176
rect 798 313824 559200 317896
rect 798 313544 559120 313824
rect 798 313008 559200 313544
rect 880 312728 559200 313008
rect 798 307840 559200 312728
rect 880 307560 559200 307840
rect 798 306752 559200 307560
rect 798 306472 559120 306752
rect 798 302672 559200 306472
rect 880 302392 559200 302672
rect 798 299680 559200 302392
rect 798 299400 559120 299680
rect 798 297504 559200 299400
rect 880 297224 559200 297504
rect 798 292608 559200 297224
rect 798 292336 559120 292608
rect 880 292328 559120 292336
rect 880 292056 559200 292328
rect 798 287168 559200 292056
rect 880 286888 559200 287168
rect 798 285536 559200 286888
rect 798 285256 559120 285536
rect 798 282000 559200 285256
rect 880 281720 559200 282000
rect 798 278464 559200 281720
rect 798 278184 559120 278464
rect 798 276832 559200 278184
rect 880 276552 559200 276832
rect 798 271664 559200 276552
rect 880 271392 559200 271664
rect 880 271384 559120 271392
rect 798 271112 559120 271384
rect 798 266496 559200 271112
rect 880 266216 559200 266496
rect 798 264320 559200 266216
rect 798 264040 559120 264320
rect 798 261328 559200 264040
rect 880 261048 559200 261328
rect 798 257248 559200 261048
rect 798 256968 559120 257248
rect 798 256160 559200 256968
rect 880 255880 559200 256160
rect 798 250992 559200 255880
rect 880 250712 559200 250992
rect 798 250176 559200 250712
rect 798 249896 559120 250176
rect 798 245824 559200 249896
rect 880 245544 559200 245824
rect 798 243104 559200 245544
rect 798 242824 559120 243104
rect 798 240656 559200 242824
rect 880 240376 559200 240656
rect 798 236032 559200 240376
rect 798 235752 559120 236032
rect 798 235488 559200 235752
rect 880 235208 559200 235488
rect 798 230320 559200 235208
rect 880 230040 559200 230320
rect 798 228960 559200 230040
rect 798 228680 559120 228960
rect 798 225152 559200 228680
rect 880 224872 559200 225152
rect 798 221888 559200 224872
rect 798 221608 559120 221888
rect 798 219984 559200 221608
rect 880 219704 559200 219984
rect 798 214816 559200 219704
rect 880 214536 559120 214816
rect 798 209648 559200 214536
rect 880 209368 559200 209648
rect 798 207744 559200 209368
rect 798 207464 559120 207744
rect 798 204480 559200 207464
rect 880 204200 559200 204480
rect 798 200672 559200 204200
rect 798 200392 559120 200672
rect 798 199312 559200 200392
rect 880 199032 559200 199312
rect 798 194144 559200 199032
rect 880 193864 559200 194144
rect 798 193600 559200 193864
rect 798 193320 559120 193600
rect 798 188976 559200 193320
rect 880 188696 559200 188976
rect 798 186528 559200 188696
rect 798 186248 559120 186528
rect 798 183808 559200 186248
rect 880 183528 559200 183808
rect 798 179456 559200 183528
rect 798 179176 559120 179456
rect 798 178640 559200 179176
rect 880 178360 559200 178640
rect 798 173472 559200 178360
rect 880 173192 559200 173472
rect 798 172384 559200 173192
rect 798 172104 559120 172384
rect 798 168304 559200 172104
rect 880 168024 559200 168304
rect 798 165312 559200 168024
rect 798 165032 559120 165312
rect 798 163136 559200 165032
rect 880 162856 559200 163136
rect 798 158240 559200 162856
rect 798 157968 559120 158240
rect 880 157960 559120 157968
rect 880 157688 559200 157960
rect 798 152800 559200 157688
rect 880 152520 559200 152800
rect 798 151168 559200 152520
rect 798 150888 559120 151168
rect 798 147632 559200 150888
rect 880 147352 559200 147632
rect 798 144096 559200 147352
rect 798 143816 559120 144096
rect 798 142464 559200 143816
rect 880 142184 559200 142464
rect 798 137296 559200 142184
rect 880 137024 559200 137296
rect 880 137016 559120 137024
rect 798 136744 559120 137016
rect 798 132128 559200 136744
rect 880 131848 559200 132128
rect 798 129952 559200 131848
rect 798 129672 559120 129952
rect 798 126960 559200 129672
rect 880 126680 559200 126960
rect 798 122880 559200 126680
rect 798 122600 559120 122880
rect 798 121792 559200 122600
rect 880 121512 559200 121792
rect 798 116624 559200 121512
rect 880 116344 559200 116624
rect 798 115808 559200 116344
rect 798 115528 559120 115808
rect 798 111456 559200 115528
rect 880 111176 559200 111456
rect 798 108736 559200 111176
rect 798 108456 559120 108736
rect 798 106288 559200 108456
rect 880 106008 559200 106288
rect 798 101664 559200 106008
rect 798 101384 559120 101664
rect 798 101120 559200 101384
rect 880 100840 559200 101120
rect 798 95952 559200 100840
rect 880 95672 559200 95952
rect 798 94592 559200 95672
rect 798 94312 559120 94592
rect 798 90784 559200 94312
rect 880 90504 559200 90784
rect 798 87520 559200 90504
rect 798 87240 559120 87520
rect 798 85616 559200 87240
rect 880 85336 559200 85616
rect 798 80448 559200 85336
rect 880 80168 559120 80448
rect 798 75280 559200 80168
rect 880 75000 559200 75280
rect 798 73376 559200 75000
rect 798 73096 559120 73376
rect 798 70112 559200 73096
rect 880 69832 559200 70112
rect 798 66304 559200 69832
rect 798 66024 559120 66304
rect 798 64944 559200 66024
rect 880 64664 559200 64944
rect 798 59776 559200 64664
rect 880 59496 559200 59776
rect 798 59232 559200 59496
rect 798 58952 559120 59232
rect 798 54608 559200 58952
rect 880 54328 559200 54608
rect 798 52160 559200 54328
rect 798 51880 559120 52160
rect 798 49440 559200 51880
rect 880 49160 559200 49440
rect 798 45088 559200 49160
rect 798 44808 559120 45088
rect 798 44272 559200 44808
rect 880 43992 559200 44272
rect 798 39104 559200 43992
rect 880 38824 559200 39104
rect 798 38016 559200 38824
rect 798 37736 559120 38016
rect 798 33936 559200 37736
rect 880 33656 559200 33936
rect 798 30944 559200 33656
rect 798 30664 559120 30944
rect 798 28768 559200 30664
rect 880 28488 559200 28768
rect 798 23872 559200 28488
rect 798 23600 559120 23872
rect 880 23592 559120 23600
rect 880 23320 559200 23592
rect 798 18432 559200 23320
rect 880 18152 559200 18432
rect 798 16800 559200 18152
rect 798 16520 559120 16800
rect 798 13264 559200 16520
rect 880 12984 559200 13264
rect 798 9728 559200 12984
rect 798 9448 559120 9728
rect 798 8096 559200 9448
rect 880 7816 559200 8096
rect 798 171 559200 7816
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 85435 2048 96288 26893
rect 96768 2048 111648 26893
rect 112128 2048 127008 26893
rect 127488 2048 142368 26893
rect 142848 2048 157728 26893
rect 158208 2048 173088 26893
rect 173568 2048 188448 26893
rect 188928 2048 203808 26893
rect 204288 2048 219168 26893
rect 219648 2048 234528 26893
rect 235008 2048 249888 26893
rect 250368 2048 265248 26893
rect 265728 2048 280608 26893
rect 281088 2048 295968 26893
rect 296448 2048 311328 26893
rect 311808 2048 326688 26893
rect 327168 2048 342048 26893
rect 342528 2048 357408 26893
rect 357888 2048 372768 26893
rect 373248 2048 388128 26893
rect 388608 2048 403488 26893
rect 403968 2048 418848 26893
rect 419328 2048 423693 26893
rect 85435 171 423693 2048
<< labels >>
rlabel metal3 s 559200 9528 560000 9648 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 559200 221688 560000 221808 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 559200 242904 560000 243024 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 559200 264120 560000 264240 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 559200 285336 560000 285456 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 559200 306552 560000 306672 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 559200 327768 560000 327888 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 343816 800 343936 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 328312 800 328432 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 312808 800 312928 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 297304 800 297424 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 559200 30744 560000 30864 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 281800 800 281920 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 266296 800 266416 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 250792 800 250912 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 235288 800 235408 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 219784 800 219904 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 204280 800 204400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 188776 800 188896 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 173272 800 173392 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 559200 51960 560000 52080 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 559200 73176 560000 73296 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 559200 94392 560000 94512 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 559200 115608 560000 115728 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 559200 136824 560000 136944 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 559200 158040 560000 158160 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 559200 179256 560000 179376 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 559200 200472 560000 200592 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 559200 23672 560000 23792 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 559200 235832 560000 235952 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 559200 257048 560000 257168 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 559200 278264 560000 278384 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 559200 299480 560000 299600 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 559200 320696 560000 320816 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 559200 341912 560000 342032 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 0 333480 800 333600 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 0 317976 800 318096 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 0 302472 800 302592 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 286968 800 287088 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 559200 44888 560000 45008 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 271464 800 271584 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 255960 800 256080 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 240456 800 240576 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 224952 800 225072 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 193944 800 194064 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 178440 800 178560 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 162936 800 163056 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 147432 800 147552 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 559200 66104 560000 66224 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 559200 87320 560000 87440 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 559200 108536 560000 108656 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 559200 129752 560000 129872 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 559200 150968 560000 151088 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 559200 172184 560000 172304 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 559200 193400 560000 193520 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 559200 214616 560000 214736 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 559200 16600 560000 16720 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 559200 228760 560000 228880 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 559200 249976 560000 250096 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 559200 271192 560000 271312 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 559200 292408 560000 292528 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 559200 313624 560000 313744 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 559200 334840 560000 334960 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 0 338648 800 338768 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 0 323144 800 323264 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 0 307640 800 307760 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 292136 800 292256 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 559200 37816 560000 37936 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 276632 800 276752 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 261128 800 261248 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 245624 800 245744 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 230120 800 230240 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 214616 800 214736 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 199112 800 199232 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 559200 59032 560000 59152 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 559200 80248 560000 80368 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 559200 101464 560000 101584 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 559200 122680 560000 122800 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 559200 143896 560000 144016 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 559200 165112 560000 165232 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 559200 186328 560000 186448 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 559200 207544 560000 207664 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 548798 0 548854 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 549902 0 549958 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 551006 0 551062 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 459374 0 459430 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 462686 0 462742 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 465998 0 466054 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 469310 0 469366 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 472622 0 472678 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 475934 0 475990 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 479246 0 479302 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 482558 0 482614 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 485870 0 485926 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 489182 0 489238 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 492494 0 492550 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 495806 0 495862 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 499118 0 499174 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 502430 0 502486 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 505742 0 505798 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 509054 0 509110 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 512366 0 512422 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 515678 0 515734 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 518990 0 519046 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 522302 0 522358 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 525614 0 525670 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 528926 0 528982 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 532238 0 532294 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 535550 0 535606 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 538862 0 538918 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 542174 0 542230 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 545486 0 545542 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 164606 0 164662 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 210974 0 211030 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 214286 0 214342 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 247406 0 247462 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 257342 0 257398 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 280526 0 280582 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 283838 0 283894 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 287150 0 287206 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 290462 0 290518 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 293774 0 293830 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 303710 0 303766 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 307022 0 307078 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 313646 0 313702 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 320270 0 320326 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 323582 0 323638 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 326894 0 326950 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 330206 0 330262 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 333518 0 333574 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 336830 0 336886 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 340142 0 340198 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 343454 0 343510 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 346766 0 346822 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 350078 0 350134 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 353390 0 353446 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 356702 0 356758 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 360014 0 360070 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 363326 0 363382 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 366638 0 366694 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 369950 0 370006 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 373262 0 373318 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 376574 0 376630 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 379886 0 379942 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 383198 0 383254 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 389822 0 389878 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 393134 0 393190 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 396446 0 396502 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 399758 0 399814 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 406382 0 406438 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 409694 0 409750 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 413006 0 413062 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 416318 0 416374 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 419630 0 419686 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 422942 0 422998 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 426254 0 426310 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 429566 0 429622 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 432878 0 432934 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 436190 0 436246 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 439502 0 439558 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 442814 0 442870 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 446126 0 446182 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 449438 0 449494 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 452750 0 452806 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 457166 0 457222 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 460478 0 460534 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 463790 0 463846 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 467102 0 467158 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 470414 0 470470 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 473726 0 473782 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 477038 0 477094 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 480350 0 480406 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 483662 0 483718 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 486974 0 487030 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 490286 0 490342 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 493598 0 493654 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 496910 0 496966 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 500222 0 500278 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 503534 0 503590 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 506846 0 506902 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 510158 0 510214 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 513470 0 513526 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 516782 0 516838 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 520094 0 520150 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 523406 0 523462 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 526718 0 526774 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 530030 0 530086 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 533342 0 533398 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 536654 0 536710 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 539966 0 540022 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 543278 0 543334 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 546590 0 546646 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 175646 0 175702 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 178958 0 179014 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 185582 0 185638 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 188894 0 188950 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 192206 0 192262 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 208766 0 208822 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 212078 0 212134 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 218702 0 218758 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 222014 0 222070 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 231950 0 232006 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 235262 0 235318 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 238574 0 238630 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 241886 0 241942 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 245198 0 245254 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 248510 0 248566 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 251822 0 251878 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 255134 0 255190 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 258446 0 258502 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 261758 0 261814 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 265070 0 265126 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 268382 0 268438 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 271694 0 271750 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 275006 0 275062 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 278318 0 278374 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 281630 0 281686 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 284942 0 284998 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 288254 0 288310 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 291566 0 291622 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 294878 0 294934 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 298190 0 298246 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 301502 0 301558 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 304814 0 304870 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 308126 0 308182 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 311438 0 311494 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 314750 0 314806 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 318062 0 318118 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 321374 0 321430 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 324686 0 324742 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 327998 0 328054 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 331310 0 331366 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 334622 0 334678 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 337934 0 337990 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 341246 0 341302 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 344558 0 344614 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 347870 0 347926 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 351182 0 351238 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 354494 0 354550 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 357806 0 357862 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 361118 0 361174 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 364430 0 364486 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 367742 0 367798 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 371054 0 371110 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 374366 0 374422 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 380990 0 381046 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 384302 0 384358 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 387614 0 387670 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 390926 0 390982 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 394238 0 394294 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 397550 0 397606 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 400862 0 400918 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 404174 0 404230 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 407486 0 407542 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 410798 0 410854 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 414110 0 414166 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 417422 0 417478 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 420734 0 420790 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 424046 0 424102 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 427358 0 427414 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 430670 0 430726 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 433982 0 434038 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 437294 0 437350 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 440606 0 440662 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 443918 0 443974 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 447230 0 447286 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 450542 0 450598 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 453854 0 453910 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 458270 0 458326 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 461582 0 461638 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 464894 0 464950 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 468206 0 468262 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 471518 0 471574 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 474830 0 474886 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 478142 0 478198 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 481454 0 481510 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 484766 0 484822 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 488078 0 488134 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 491390 0 491446 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 494702 0 494758 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 498014 0 498070 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 501326 0 501382 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 504638 0 504694 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 507950 0 508006 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 511262 0 511318 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 514574 0 514630 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 517886 0 517942 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 521198 0 521254 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 524510 0 524566 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 527822 0 527878 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 531134 0 531190 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 534446 0 534502 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 537758 0 537814 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 541070 0 541126 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 544382 0 544438 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 547694 0 547750 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 193310 0 193366 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 252926 0 252982 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 262862 0 262918 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 272798 0 272854 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 286046 0 286102 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 289358 0 289414 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 309230 0 309286 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 319166 0 319222 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 332414 0 332470 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 335726 0 335782 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 342350 0 342406 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 345662 0 345718 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 348974 0 349030 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 355598 0 355654 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 358910 0 358966 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 362222 0 362278 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 368846 0 368902 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 372158 0 372214 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 375470 0 375526 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 378782 0 378838 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 382094 0 382150 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 385406 0 385462 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 392030 0 392086 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 395342 0 395398 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 398654 0 398710 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 401966 0 402022 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 405278 0 405334 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 408590 0 408646 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 415214 0 415270 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 418526 0 418582 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 421838 0 421894 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 425150 0 425206 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 428462 0 428518 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 431774 0 431830 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 435086 0 435142 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 438398 0 438454 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 441710 0 441766 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 445022 0 445078 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 448334 0 448390 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 451646 0 451702 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 454958 0 455014 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 552110 0 552166 800 6 user_clock2
port 502 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 504 nsew ground bidirectional
rlabel metal2 s 7838 0 7894 800 6 wb_clk_i
port 505 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb_rst_i
port 506 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_ack_o
port 507 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[0]
port 508 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_adr_i[10]
port 509 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 wbs_adr_i[11]
port 510 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wbs_adr_i[12]
port 511 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_adr_i[13]
port 512 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 wbs_adr_i[14]
port 513 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[15]
port 514 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_adr_i[16]
port 515 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_adr_i[17]
port 516 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_adr_i[18]
port 517 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_adr_i[19]
port 518 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[1]
port 519 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 wbs_adr_i[20]
port 520 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wbs_adr_i[21]
port 521 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 wbs_adr_i[22]
port 522 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 wbs_adr_i[23]
port 523 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_adr_i[24]
port 524 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 wbs_adr_i[25]
port 525 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_adr_i[26]
port 526 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wbs_adr_i[27]
port 527 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_adr_i[28]
port 528 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_adr_i[29]
port 529 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_adr_i[2]
port 530 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 wbs_adr_i[30]
port 531 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 wbs_adr_i[31]
port 532 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[3]
port 533 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_adr_i[4]
port 534 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[5]
port 535 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_adr_i[6]
port 536 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[7]
port 537 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_adr_i[8]
port 538 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[9]
port 539 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_cyc_i
port 540 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[0]
port 541 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[10]
port 542 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_i[11]
port 543 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[12]
port 544 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_i[13]
port 545 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[14]
port 546 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_i[15]
port 547 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 wbs_dat_i[16]
port 548 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 wbs_dat_i[17]
port 549 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_i[18]
port 550 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 wbs_dat_i[19]
port 551 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[1]
port 552 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_dat_i[20]
port 553 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 wbs_dat_i[21]
port 554 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 wbs_dat_i[22]
port 555 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_dat_i[23]
port 556 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wbs_dat_i[24]
port 557 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_i[25]
port 558 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[26]
port 559 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 wbs_dat_i[27]
port 560 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 wbs_dat_i[28]
port 561 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_i[29]
port 562 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[2]
port 563 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 wbs_dat_i[30]
port 564 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[31]
port 565 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[3]
port 566 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[4]
port 567 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[5]
port 568 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[6]
port 569 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_i[7]
port 570 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_i[8]
port 571 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_i[9]
port 572 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[0]
port 573 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_o[10]
port 574 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 wbs_dat_o[11]
port 575 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_o[12]
port 576 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[13]
port 577 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_o[14]
port 578 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 wbs_dat_o[15]
port 579 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_o[16]
port 580 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 wbs_dat_o[17]
port 581 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_o[18]
port 582 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 wbs_dat_o[19]
port 583 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[1]
port 584 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 wbs_dat_o[20]
port 585 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 wbs_dat_o[21]
port 586 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 wbs_dat_o[22]
port 587 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 wbs_dat_o[23]
port 588 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 wbs_dat_o[24]
port 589 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 wbs_dat_o[25]
port 590 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 wbs_dat_o[26]
port 591 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_o[27]
port 592 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 wbs_dat_o[28]
port 593 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 wbs_dat_o[29]
port 594 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[2]
port 595 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 wbs_dat_o[30]
port 596 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 wbs_dat_o[31]
port 597 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_o[3]
port 598 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[4]
port 599 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_o[5]
port 600 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[6]
port 601 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_o[7]
port 602 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[8]
port 603 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_o[9]
port 604 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_stb_i
port 609 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_we_i
port 610 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68017250
string GDS_FILE /home/ucass/Work/DNN_ACC_IITGN/openlane/user_proj_mac/runs/23_09_23_01_27/results/signoff/user_proj_mac.magic.gds
string GDS_START 1057110
<< end >>

